-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_45_load_0_req_0 : boolean;
  signal ptr_deref_45_load_0_ack_0 : boolean;
  signal ptr_deref_45_load_0_req_1 : boolean;
  signal ptr_deref_45_load_0_ack_1 : boolean;
  signal ptr_deref_57_load_0_req_0 : boolean;
  signal ptr_deref_57_load_0_ack_0 : boolean;
  signal ptr_deref_57_load_0_req_1 : boolean;
  signal ptr_deref_57_load_0_ack_1 : boolean;
  signal type_cast_171_inst_req_0 : boolean;
  signal type_cast_171_inst_ack_0 : boolean;
  signal type_cast_171_inst_req_1 : boolean;
  signal type_cast_171_inst_ack_1 : boolean;
  signal ptr_deref_69_load_0_req_0 : boolean;
  signal ptr_deref_69_load_0_ack_0 : boolean;
  signal ptr_deref_69_load_0_req_1 : boolean;
  signal ptr_deref_69_load_0_ack_1 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal if_stmt_98_branch_req_0 : boolean;
  signal if_stmt_98_branch_ack_1 : boolean;
  signal if_stmt_98_branch_ack_0 : boolean;
  signal type_cast_117_inst_req_0 : boolean;
  signal type_cast_117_inst_ack_0 : boolean;
  signal type_cast_117_inst_req_1 : boolean;
  signal type_cast_117_inst_ack_1 : boolean;
  signal array_obj_ref_152_index_offset_req_0 : boolean;
  signal array_obj_ref_152_index_offset_ack_0 : boolean;
  signal array_obj_ref_152_index_offset_req_1 : boolean;
  signal array_obj_ref_152_index_offset_ack_1 : boolean;
  signal addr_of_153_final_reg_req_0 : boolean;
  signal addr_of_153_final_reg_ack_0 : boolean;
  signal addr_of_153_final_reg_req_1 : boolean;
  signal addr_of_153_final_reg_ack_1 : boolean;
  signal ptr_deref_157_load_0_req_0 : boolean;
  signal ptr_deref_157_load_0_ack_0 : boolean;
  signal ptr_deref_157_load_0_req_1 : boolean;
  signal ptr_deref_157_load_0_ack_1 : boolean;
  signal type_cast_161_inst_req_0 : boolean;
  signal type_cast_161_inst_ack_0 : boolean;
  signal type_cast_161_inst_req_1 : boolean;
  signal type_cast_161_inst_ack_1 : boolean;
  signal type_cast_181_inst_req_0 : boolean;
  signal type_cast_181_inst_ack_0 : boolean;
  signal type_cast_181_inst_req_1 : boolean;
  signal type_cast_181_inst_ack_1 : boolean;
  signal type_cast_191_inst_req_0 : boolean;
  signal type_cast_191_inst_ack_0 : boolean;
  signal type_cast_191_inst_req_1 : boolean;
  signal type_cast_191_inst_ack_1 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal type_cast_221_inst_req_0 : boolean;
  signal type_cast_221_inst_ack_0 : boolean;
  signal type_cast_221_inst_req_1 : boolean;
  signal type_cast_221_inst_ack_1 : boolean;
  signal type_cast_231_inst_req_0 : boolean;
  signal type_cast_231_inst_ack_0 : boolean;
  signal type_cast_231_inst_req_1 : boolean;
  signal type_cast_231_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_248_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_248_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_248_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_248_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_251_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_251_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_251_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_251_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_254_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_254_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_254_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_254_inst_ack_1 : boolean;
  signal if_stmt_268_branch_req_0 : boolean;
  signal if_stmt_268_branch_ack_1 : boolean;
  signal if_stmt_268_branch_ack_0 : boolean;
  signal phi_stmt_140_req_0 : boolean;
  signal type_cast_146_inst_req_0 : boolean;
  signal type_cast_146_inst_ack_0 : boolean;
  signal type_cast_146_inst_req_1 : boolean;
  signal type_cast_146_inst_ack_1 : boolean;
  signal phi_stmt_140_req_1 : boolean;
  signal phi_stmt_140_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(68);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	9 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_34/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/branch_block_stmt_34__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Update/cr
      -- 
    rr_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_45_load_0_req_0); -- 
    cr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_45_load_0_req_1); -- 
    rr_139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_57_load_0_req_0); -- 
    cr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_57_load_0_req_1); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_69_load_0_req_0); -- 
    cr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_69_load_0_req_1); -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_83_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Sample/word_access_start/word_0/ra
      -- 
    ra_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_45_load_0_ack_0, ack => sendOutput_CP_26_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/ptr_deref_45_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/ptr_deref_45_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/ptr_deref_45_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_45_Update/ptr_deref_45_Merge/merge_ack
      -- 
    ca_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_45_load_0_ack_1, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Sample/word_access_start/word_0/ra
      -- 
    ra_140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_57_load_0_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/ptr_deref_57_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/ptr_deref_57_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/ptr_deref_57_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_57_Update/ptr_deref_57_Merge/merge_ack
      -- 
    ca_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_57_load_0_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Sample/word_access_start/word_0/ra
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_69_load_0_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/ptr_deref_69_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/ptr_deref_69_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/ptr_deref_69_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/ptr_deref_69_Update/ptr_deref_69_Merge/merge_ack
      -- 
    ca_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_69_load_0_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Sample/rr
      -- 
    rr_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(7), ack => type_cast_83_inst_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(6) & sendOutput_CP_26_elements(2) & sendOutput_CP_26_elements(4);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Sample/ra
      -- 
    ra_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => sendOutput_CP_26_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (13) 
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97__exit__
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98__entry__
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/$exit
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_42_to_assign_stmt_97/type_cast_83_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_34/R_cmp77_99_place
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/if_stmt_98_else_link/$entry
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => sendOutput_CP_26_elements(9)); -- 
    branch_req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(9), ack => if_stmt_98_branch_req_0); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	68 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_34/if_stmt_98_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_34/if_stmt_98_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_34/entry_forx_xend
      -- CP-element group 10: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_98_branch_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (18) 
      -- CP-element group 11: 	 branch_block_stmt_34/merge_stmt_104__exit__
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137__entry__
      -- CP-element group 11: 	 branch_block_stmt_34/if_stmt_98_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/if_stmt_98_else_link/else_choice_transition
      -- CP-element group 11: 	 branch_block_stmt_34/entry_bbx_xnph
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/$entry
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_update_start_
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_34/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_34/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/merge_stmt_104_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_34/merge_stmt_104_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_34/merge_stmt_104_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/merge_stmt_104_PhiAck/dummy
      -- 
    else_choice_transition_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_98_branch_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_117_inst_req_0); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_117_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_117_inst_ack_0, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  place  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	62 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137__exit__
      -- CP-element group 13: 	 branch_block_stmt_34/bbx_xnph_forx_xbody
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/$exit
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_109_to_assign_stmt_137/type_cast_117_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/phi_stmt_140/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/$entry
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_117_inst_ack_1, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	59 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_sample_complete
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Sample/ack
      -- 
    ack_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_152_index_offset_ack_0, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	67 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (11) 
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Update/ack
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_request/$entry
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_request/req
      -- 
    ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_152_index_offset_ack_1, ack => sendOutput_CP_26_elements(15)); -- 
    req_299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => addr_of_153_final_reg_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_request/$exit
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_request/ack
      -- 
    ack_300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_153_final_reg_ack_0, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (24) 
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_complete/ack
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_word_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_address_resized
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_addr_resize/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_addr_resize/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_addr_resize/base_resize_req
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_addr_resize/base_resize_ack
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_word_addrgen/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_word_addrgen/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_word_addrgen/root_register_req
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_word_addrgen/root_register_ack
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/word_access_start/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/word_access_start/word_0/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/word_access_start/word_0/rr
      -- 
    ack_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_153_final_reg_ack_1, ack => sendOutput_CP_26_elements(17)); -- 
    rr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(17), ack => ptr_deref_157_load_0_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/word_access_start/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Sample/word_access_start/word_0/ra
      -- 
    ra_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_157_load_0_ack_0, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	67 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	28 
    -- CP-element group 19: 	30 
    -- CP-element group 19: 	32 
    -- CP-element group 19: 	34 
    -- CP-element group 19: 	24 
    -- CP-element group 19:  members (33) 
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/word_access_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/ptr_deref_157_Merge/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/ptr_deref_157_Merge/$exit
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/ptr_deref_157_Merge/merge_req
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/ptr_deref_157_Merge/merge_ack
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Sample/rr
      -- 
    ca_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_157_load_0_ack_1, ack => sendOutput_CP_26_elements(19)); -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_171_inst_req_0); -- 
    rr_405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_191_inst_req_0); -- 
    rr_419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_201_inst_req_0); -- 
    rr_433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_211_inst_req_0); -- 
    rr_447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_221_inst_req_0); -- 
    rr_461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_231_inst_req_0); -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_161_inst_req_0); -- 
    rr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_181_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Sample/ra
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_161_inst_ack_0, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	67 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Update/ca
      -- 
    ca_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_161_inst_ack_1, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Sample/$exit
      -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_171_inst_ack_0, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	67 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	53 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_update_completed_
      -- 
    ca_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_171_inst_ack_1, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Sample/ra
      -- 
    ra_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_0, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	67 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Update/ca
      -- 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_1, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Sample/ra
      -- 
    ra_406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_191_inst_ack_0, ack => sendOutput_CP_26_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	67 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	47 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Update/ca
      -- 
    ca_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_191_inst_ack_1, ack => sendOutput_CP_26_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Sample/ra
      -- 
    ra_420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	44 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Update/ca
      -- 
    ca_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => sendOutput_CP_26_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	19 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Sample/ra
      -- 
    ra_434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	67 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	41 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Update/ca
      -- 
    ca_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	19 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Sample/ra
      -- 
    ra_448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_221_inst_ack_0, ack => sendOutput_CP_26_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	67 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Update/ca
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_221_inst_ack_1, ack => sendOutput_CP_26_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Sample/ra
      -- 
    ra_462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_231_inst_ack_0, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	67 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Sample/req
      -- 
    ca_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_231_inst_ack_1, ack => sendOutput_CP_26_elements(35)); -- 
    req_475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_233_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_update_start_
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Update/req
      -- 
    ack_476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_233_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_233_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_233_Update/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_233_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Sample/req
      -- 
    req_489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_236_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(33) & sendOutput_CP_26_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_update_start_
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Update/req
      -- 
    ack_490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_236_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_236_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_236_Update/ack
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_236_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	31 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Sample/req
      -- 
    req_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_239_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(31) & sendOutput_CP_26_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_update_start_
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Update/req
      -- 
    ack_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_239_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_239_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_239_Update/ack
      -- 
    ack_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_239_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Sample/req
      -- 
    req_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_242_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(29) & sendOutput_CP_26_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_update_start_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Update/req
      -- 
    ack_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_242_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_242_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_242_Update/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_242_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	27 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Sample/req
      -- 
    req_531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_245_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(27) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_update_start_
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Update/req
      -- 
    ack_532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_245_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_245_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_245_Update/ack
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_245_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Sample/req
      -- 
    req_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => WPIPE_zeropad_output_pipe_248_inst_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(25) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_update_start_
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Update/req
      -- 
    ack_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_248_inst_ack_0, ack => sendOutput_CP_26_elements(51)); -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(51), ack => WPIPE_zeropad_output_pipe_248_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_248_Update/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_248_inst_ack_1, ack => sendOutput_CP_26_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	23 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Sample/req
      -- 
    req_559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => WPIPE_zeropad_output_pipe_251_inst_req_0); -- 
    sendOutput_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(52) & sendOutput_CP_26_elements(23);
      gj_sendOutput_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_update_start_
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Update/req
      -- 
    ack_560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_251_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(54), ack => WPIPE_zeropad_output_pipe_251_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_251_Update/ack
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_251_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Sample/req
      -- 
    req_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => WPIPE_zeropad_output_pipe_254_inst_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(21) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_update_start_
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Update/req
      -- 
    ack_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_254_inst_ack_0, ack => sendOutput_CP_26_elements(57)); -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(57), ack => WPIPE_zeropad_output_pipe_254_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/WPIPE_zeropad_output_pipe_254_Update/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_254_inst_ack_1, ack => sendOutput_CP_26_elements(58)); -- 
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267__exit__
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268__entry__
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/$exit
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_34/R_exitcond9_269_place
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/if_stmt_268_else_link/$entry
      -- 
    branch_req_587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(59), ack => if_stmt_268_branch_req_0); -- 
    sendOutput_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(14) & sendOutput_CP_26_elements(58);
      gj_sendOutput_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  merge  transition  place  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_34/merge_stmt_274__exit__
      -- CP-element group 60: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend
      -- CP-element group 60: 	 branch_block_stmt_34/if_stmt_268_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/if_stmt_268_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 60: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/merge_stmt_274_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_34/merge_stmt_274_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_34/merge_stmt_274_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/merge_stmt_274_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_268_branch_ack_1, ack => sendOutput_CP_26_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	64 
    -- CP-element group 61:  members (12) 
      -- CP-element group 61: 	 branch_block_stmt_34/if_stmt_268_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/if_stmt_268_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Update/cr
      -- 
    else_choice_transition_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_268_branch_ack_0, ack => sendOutput_CP_26_elements(61)); -- 
    rr_640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_146_inst_req_0); -- 
    cr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_146_inst_req_1); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	13 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/phi_stmt_140/$exit
      -- CP-element group 62: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_144_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_34/bbx_xnph_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_req
      -- 
    phi_stmt_140_req_621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_140_req_621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(62), ack => phi_stmt_140_req_0); -- 
    -- Element group sendOutput_CP_26_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(13), ack => sendOutput_CP_26_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Sample/ra
      -- 
    ra_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_0, ack => sendOutput_CP_26_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	61 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/Update/ca
      -- 
    ca_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_1, ack => sendOutput_CP_26_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_sources/type_cast_146/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_140/phi_stmt_140_req
      -- 
    phi_stmt_140_req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_140_req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(65), ack => phi_stmt_140_req_1); -- 
    sendOutput_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(63) & sendOutput_CP_26_elements(64);
      gj_sendOutput_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_34/merge_stmt_139_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_34/merge_stmt_139_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(66) <= OrReduce(sendOutput_CP_26_elements(62) & sendOutput_CP_26_elements(65));
    -- CP-element group 67:  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	21 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	27 
    -- CP-element group 67: 	29 
    -- CP-element group 67: 	31 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	35 
    -- CP-element group 67: 	19 
    -- CP-element group 67: 	23 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	14 
    -- CP-element group 67: 	15 
    -- CP-element group 67:  members (53) 
      -- CP-element group 67: 	 branch_block_stmt_34/merge_stmt_139__exit__
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267__entry__
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_resized_1
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_scaled_1
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_computed_1
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_resize_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_resize_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_resize_1/index_resize_req
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_resize_1/index_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_scale_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_scale_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_scale_1/scale_rename_req
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_index_scale_1/scale_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_update_start
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/array_obj_ref_152_final_index_sum_regn_Update/req
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/addr_of_153_complete/req
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/word_access_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/word_access_complete/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/ptr_deref_157_Update/word_access_complete/word_0/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_161_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_171_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_181_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_191_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_201_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_211_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_221_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_update_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_154_to_assign_stmt_267/type_cast_231_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_34/merge_stmt_139_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_34/merge_stmt_139_PhiAck/phi_stmt_140_ack
      -- 
    phi_stmt_140_ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_140_ack_0, ack => sendOutput_CP_26_elements(67)); -- 
    cr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_171_inst_req_1); -- 
    req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_152_index_offset_req_0); -- 
    req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_152_index_offset_req_1); -- 
    req_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => addr_of_153_final_reg_req_1); -- 
    cr_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => ptr_deref_157_load_0_req_1); -- 
    cr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_161_inst_req_1); -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_181_inst_req_1); -- 
    cr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_191_inst_req_1); -- 
    cr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_201_inst_req_1); -- 
    cr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_211_inst_req_1); -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_221_inst_req_1); -- 
    cr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_231_inst_req_1); -- 
    -- CP-element group 68:  merge  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	10 
    -- CP-element group 68: 	60 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_34/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/branch_block_stmt_34__exit__
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_276__exit__
      -- CP-element group 68: 	 branch_block_stmt_34/return__
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_278__exit__
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_276_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_276_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_276_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_276_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_34/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_34/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_278_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_278_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_278_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/merge_stmt_278_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(68) <= OrReduce(sendOutput_CP_26_elements(10) & sendOutput_CP_26_elements(60));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_151_resized : std_logic_vector(13 downto 0);
    signal R_indvar_151_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_152_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_152_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_152_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_152_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_152_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_152_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_154 : std_logic_vector(31 downto 0);
    signal cmp77_97 : std_logic_vector(0 downto 0);
    signal conv14_162 : std_logic_vector(7 downto 0);
    signal conv20_172 : std_logic_vector(7 downto 0);
    signal conv26_182 : std_logic_vector(7 downto 0);
    signal conv32_192 : std_logic_vector(7 downto 0);
    signal conv38_202 : std_logic_vector(7 downto 0);
    signal conv44_212 : std_logic_vector(7 downto 0);
    signal conv50_222 : std_logic_vector(7 downto 0);
    signal conv56_232 : std_logic_vector(7 downto 0);
    signal conv_84 : std_logic_vector(63 downto 0);
    signal exitcond9_267 : std_logic_vector(0 downto 0);
    signal iNsTr_0_42 : std_logic_vector(31 downto 0);
    signal iNsTr_1_54 : std_logic_vector(31 downto 0);
    signal iNsTr_2_66 : std_logic_vector(31 downto 0);
    signal indvar_140 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_262 : std_logic_vector(63 downto 0);
    signal mul3_80 : std_logic_vector(31 downto 0);
    signal mul_75 : std_logic_vector(31 downto 0);
    signal ptr_deref_157_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_157_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_157_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_157_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_157_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_45_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_45_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_45_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_45_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_45_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_57_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_57_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_57_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_57_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_57_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_69_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_69_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_69_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_69_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_69_word_offset_0 : std_logic_vector(6 downto 0);
    signal shr17_168 : std_logic_vector(63 downto 0);
    signal shr23_178 : std_logic_vector(63 downto 0);
    signal shr29_188 : std_logic_vector(63 downto 0);
    signal shr35_198 : std_logic_vector(63 downto 0);
    signal shr41_208 : std_logic_vector(63 downto 0);
    signal shr47_218 : std_logic_vector(63 downto 0);
    signal shr53_228 : std_logic_vector(63 downto 0);
    signal shr76x_xmask_90 : std_logic_vector(63 downto 0);
    signal tmp11_158 : std_logic_vector(63 downto 0);
    signal tmp1_58 : std_logic_vector(31 downto 0);
    signal tmp2_70 : std_logic_vector(31 downto 0);
    signal tmp3_109 : std_logic_vector(31 downto 0);
    signal tmp4_114 : std_logic_vector(31 downto 0);
    signal tmp5_118 : std_logic_vector(63 downto 0);
    signal tmp6_124 : std_logic_vector(63 downto 0);
    signal tmp7_130 : std_logic_vector(0 downto 0);
    signal tmp_46 : std_logic_vector(31 downto 0);
    signal type_cast_122_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_135_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_144_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_146_wire : std_logic_vector(63 downto 0);
    signal type_cast_166_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_176_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_186_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_196_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_206_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_216_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_226_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_260_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_88_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(63 downto 0);
    signal umax8_137 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_152_constant_part_of_offset <= "00000000000000";
    array_obj_ref_152_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_152_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_152_resized_base_address <= "00000000000000";
    iNsTr_0_42 <= "00000000000000000000000000000011";
    iNsTr_1_54 <= "00000000000000000000000000000100";
    iNsTr_2_66 <= "00000000000000000000000000000101";
    ptr_deref_157_word_offset_0 <= "00000000000000";
    ptr_deref_45_word_offset_0 <= "0000000";
    ptr_deref_57_word_offset_0 <= "0000000";
    ptr_deref_69_word_offset_0 <= "0000000";
    type_cast_122_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_128_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_135_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_144_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_166_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_176_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_186_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_196_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_216_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_226_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_260_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_88_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_94_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_140: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_144_wire_constant & type_cast_146_wire;
      req <= phi_stmt_140_req_0 & phi_stmt_140_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_140",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_140_ack_0,
          idata => idata,
          odata => indvar_140,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_140
    -- flow-through select operator MUX_136_inst
    umax8_137 <= tmp6_124 when (tmp7_130(0) /=  '0') else type_cast_135_wire_constant;
    addr_of_153_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_153_final_reg_req_0;
      addr_of_153_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_153_final_reg_req_1;
      addr_of_153_final_reg_ack_1<= rack(0);
      addr_of_153_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_153_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_152_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_154,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_117_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_117_inst_req_0;
      type_cast_117_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_117_inst_req_1;
      type_cast_117_inst_ack_1<= rack(0);
      type_cast_117_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_117_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_146_inst_req_0;
      type_cast_146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_146_inst_req_1;
      type_cast_146_inst_ack_1<= rack(0);
      type_cast_146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_146_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_161_inst_req_0;
      type_cast_161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_161_inst_req_1;
      type_cast_161_inst_ack_1<= rack(0);
      type_cast_161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_171_inst_req_0;
      type_cast_171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_171_inst_req_1;
      type_cast_171_inst_ack_1<= rack(0);
      type_cast_171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_181_inst_req_0;
      type_cast_181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_181_inst_req_1;
      type_cast_181_inst_ack_1<= rack(0);
      type_cast_181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_191_inst_req_0;
      type_cast_191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_191_inst_req_1;
      type_cast_191_inst_ack_1<= rack(0);
      type_cast_191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_192,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_221_inst_req_0;
      type_cast_221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_221_inst_req_1;
      type_cast_221_inst_ack_1<= rack(0);
      type_cast_221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_231_inst_req_0;
      type_cast_231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_231_inst_req_1;
      type_cast_231_inst_ack_1<= rack(0);
      type_cast_231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr53_228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul3_80,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_84,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_152_index_1_rename
    process(R_indvar_151_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_151_resized;
      ov(13 downto 0) := iv;
      R_indvar_151_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_152_index_1_resize
    process(indvar_140) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_140;
      ov := iv(13 downto 0);
      R_indvar_151_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_152_root_address_inst
    process(array_obj_ref_152_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_152_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_152_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_addr_0
    process(ptr_deref_157_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_157_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_157_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_base_resize
    process(arrayidx_154) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_154;
      ov := iv(13 downto 0);
      ptr_deref_157_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_gather_scatter
    process(ptr_deref_157_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_157_data_0;
      ov(63 downto 0) := iv;
      tmp11_158 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_root_address_inst
    process(ptr_deref_157_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_157_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_157_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_45_addr_0
    process(ptr_deref_45_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_45_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_45_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_45_base_resize
    process(iNsTr_0_42) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_42;
      ov := iv(6 downto 0);
      ptr_deref_45_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_45_gather_scatter
    process(ptr_deref_45_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_45_data_0;
      ov(31 downto 0) := iv;
      tmp_46 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_45_root_address_inst
    process(ptr_deref_45_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_45_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_45_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_57_addr_0
    process(ptr_deref_57_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_57_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_57_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_57_base_resize
    process(iNsTr_1_54) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_54;
      ov := iv(6 downto 0);
      ptr_deref_57_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_57_gather_scatter
    process(ptr_deref_57_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_57_data_0;
      ov(31 downto 0) := iv;
      tmp1_58 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_57_root_address_inst
    process(ptr_deref_57_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_57_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_57_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_69_addr_0
    process(ptr_deref_69_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_69_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_69_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_69_base_resize
    process(iNsTr_2_66) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_66;
      ov := iv(6 downto 0);
      ptr_deref_69_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_69_gather_scatter
    process(ptr_deref_69_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_69_data_0;
      ov(31 downto 0) := iv;
      tmp2_70 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_69_root_address_inst
    process(ptr_deref_69_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_69_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_69_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_268_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_267;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_268_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_268_branch_req_0,
          ack0 => if_stmt_268_branch_ack_0,
          ack1 => if_stmt_268_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_98_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_97;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_98_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_98_branch_req_0,
          ack0 => if_stmt_98_branch_ack_0,
          ack1 => if_stmt_98_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_261_inst
    process(indvar_140) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_140, type_cast_260_wire_constant, tmp_var);
      indvarx_xnext_262 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_89_inst
    process(conv_84) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv_84, type_cast_88_wire_constant, tmp_var);
      shr76x_xmask_90 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_266_inst
    process(indvarx_xnext_262, umax8_137) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_262, umax8_137, tmp_var);
      exitcond9_267 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_95_inst
    process(shr76x_xmask_90) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr76x_xmask_90, type_cast_94_wire_constant, tmp_var);
      cmp77_97 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_123_inst
    process(tmp5_118) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_118, type_cast_122_wire_constant, tmp_var);
      tmp6_124 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_167_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_166_wire_constant, tmp_var);
      shr17_168 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_177_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_176_wire_constant, tmp_var);
      shr23_178 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_187_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_186_wire_constant, tmp_var);
      shr29_188 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_197_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_196_wire_constant, tmp_var);
      shr35_198 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_207_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_206_wire_constant, tmp_var);
      shr41_208 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_217_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_216_wire_constant, tmp_var);
      shr47_218 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_227_inst
    process(tmp11_158) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_158, type_cast_226_wire_constant, tmp_var);
      shr53_228 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_108_inst
    process(tmp1_58, tmp_46) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_58, tmp_46, tmp_var);
      tmp3_109 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_113_inst
    process(tmp3_109, tmp2_70) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_109, tmp2_70, tmp_var);
      tmp4_114 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_74_inst
    process(tmp1_58, tmp_46) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_58, tmp_46, tmp_var);
      mul_75 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_79_inst
    process(mul_75, tmp2_70) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_75, tmp2_70, tmp_var);
      mul3_80 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_129_inst
    process(tmp6_124) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp6_124, type_cast_128_wire_constant, tmp_var);
      tmp7_130 <= tmp_var; --
    end process;
    -- shared split operator group (17) : array_obj_ref_152_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_151_scaled;
      array_obj_ref_152_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_152_index_offset_req_0;
      array_obj_ref_152_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_152_index_offset_req_1;
      array_obj_ref_152_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : ptr_deref_157_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_157_load_0_req_0;
      ptr_deref_157_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_157_load_0_req_1;
      ptr_deref_157_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_157_word_address_0;
      ptr_deref_157_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_45_load_0 ptr_deref_57_load_0 ptr_deref_69_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_45_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_57_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_69_load_0_req_0;
      ptr_deref_45_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_57_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_69_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_45_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_57_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_69_load_0_req_1;
      ptr_deref_45_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_57_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_69_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_45_word_address_0 & ptr_deref_57_word_address_0 & ptr_deref_69_word_address_0;
      ptr_deref_45_data_0 <= data_out(95 downto 64);
      ptr_deref_57_data_0 <= data_out(63 downto 32);
      ptr_deref_69_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(6 downto 0),
          mtag => memory_space_4_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_233_inst WPIPE_zeropad_output_pipe_236_inst WPIPE_zeropad_output_pipe_239_inst WPIPE_zeropad_output_pipe_242_inst WPIPE_zeropad_output_pipe_245_inst WPIPE_zeropad_output_pipe_248_inst WPIPE_zeropad_output_pipe_251_inst WPIPE_zeropad_output_pipe_254_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_233_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_236_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_239_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_242_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_245_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_248_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_251_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_254_inst_req_0;
      WPIPE_zeropad_output_pipe_233_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_236_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_239_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_242_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_245_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_248_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_251_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_254_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_233_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_236_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_239_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_242_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_245_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_248_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_251_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_254_inst_req_1;
      WPIPE_zeropad_output_pipe_233_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_236_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_239_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_242_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_245_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_248_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_251_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_254_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv56_232 & conv50_222 & conv44_212 & conv38_202 & conv32_192 & conv26_182 & conv20_172 & conv14_162;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_684_start: Boolean;
  signal testConfigure_CP_684_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_615_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_296_inst_ack_0 : boolean;
  signal ptr_deref_744_store_0_req_1 : boolean;
  signal type_cast_369_inst_req_0 : boolean;
  signal array_obj_ref_607_index_offset_req_1 : boolean;
  signal type_cast_300_inst_ack_1 : boolean;
  signal type_cast_539_inst_ack_0 : boolean;
  signal if_stmt_338_branch_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_ack_1 : boolean;
  signal type_cast_615_inst_ack_1 : boolean;
  signal if_stmt_338_branch_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_696_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_611_inst_req_0 : boolean;
  signal type_cast_664_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_714_inst_req_1 : boolean;
  signal ptr_deref_525_load_0_req_1 : boolean;
  signal type_cast_369_inst_req_1 : boolean;
  signal type_cast_369_inst_ack_1 : boolean;
  signal array_obj_ref_607_index_offset_ack_1 : boolean;
  signal type_cast_317_inst_req_0 : boolean;
  signal type_cast_664_inst_req_0 : boolean;
  signal type_cast_369_inst_ack_0 : boolean;
  signal ptr_deref_525_load_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_296_inst_req_0 : boolean;
  signal type_cast_300_inst_ack_0 : boolean;
  signal ptr_deref_525_load_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_624_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_624_inst_ack_0 : boolean;
  signal if_stmt_553_branch_req_0 : boolean;
  signal type_cast_300_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_714_inst_ack_0 : boolean;
  signal type_cast_300_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_678_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_696_inst_req_0 : boolean;
  signal type_cast_539_inst_req_1 : boolean;
  signal type_cast_682_inst_req_0 : boolean;
  signal ptr_deref_309_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_732_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_714_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_624_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_624_inst_ack_1 : boolean;
  signal if_stmt_553_branch_ack_1 : boolean;
  signal type_cast_682_inst_ack_0 : boolean;
  signal ptr_deref_309_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_req_0 : boolean;
  signal ptr_deref_291_store_0_ack_1 : boolean;
  signal type_cast_700_inst_ack_0 : boolean;
  signal type_cast_718_inst_req_0 : boolean;
  signal ptr_deref_291_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_678_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_732_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_732_inst_ack_0 : boolean;
  signal type_cast_682_inst_req_1 : boolean;
  signal ptr_deref_309_store_0_ack_1 : boolean;
  signal type_cast_628_inst_req_1 : boolean;
  signal type_cast_682_inst_ack_1 : boolean;
  signal ptr_deref_525_load_0_ack_1 : boolean;
  signal type_cast_736_inst_req_0 : boolean;
  signal type_cast_664_inst_ack_1 : boolean;
  signal type_cast_317_inst_ack_1 : boolean;
  signal type_cast_317_inst_req_1 : boolean;
  signal ptr_deref_326_store_0_ack_1 : boolean;
  signal ptr_deref_744_store_0_req_0 : boolean;
  signal ptr_deref_291_store_0_ack_0 : boolean;
  signal type_cast_718_inst_ack_0 : boolean;
  signal ptr_deref_291_store_0_req_0 : boolean;
  signal type_cast_664_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_732_inst_ack_1 : boolean;
  signal array_obj_ref_607_index_offset_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_ack_0 : boolean;
  signal ptr_deref_309_store_0_req_1 : boolean;
  signal addr_of_608_final_reg_req_0 : boolean;
  signal addr_of_608_final_reg_ack_0 : boolean;
  signal array_obj_ref_607_index_offset_ack_0 : boolean;
  signal type_cast_539_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_678_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_678_inst_req_0 : boolean;
  signal type_cast_736_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_296_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_714_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_296_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_req_1 : boolean;
  signal type_cast_615_inst_req_1 : boolean;
  signal if_stmt_553_branch_ack_0 : boolean;
  signal type_cast_700_inst_req_0 : boolean;
  signal addr_of_608_final_reg_req_1 : boolean;
  signal addr_of_608_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_611_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_696_inst_ack_1 : boolean;
  signal if_stmt_338_branch_req_0 : boolean;
  signal type_cast_539_inst_req_0 : boolean;
  signal ptr_deref_326_store_0_req_0 : boolean;
  signal type_cast_317_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_req_1 : boolean;
  signal ptr_deref_326_store_0_req_1 : boolean;
  signal ptr_deref_326_store_0_ack_0 : boolean;
  signal type_cast_615_inst_ack_0 : boolean;
  signal ptr_deref_744_store_0_ack_0 : boolean;
  signal ptr_deref_744_store_0_ack_1 : boolean;
  signal type_cast_628_inst_req_0 : boolean;
  signal type_cast_628_inst_ack_0 : boolean;
  signal array_obj_ref_375_index_offset_req_0 : boolean;
  signal array_obj_ref_375_index_offset_ack_0 : boolean;
  signal array_obj_ref_375_index_offset_req_1 : boolean;
  signal array_obj_ref_375_index_offset_ack_1 : boolean;
  signal addr_of_376_final_reg_req_0 : boolean;
  signal addr_of_376_final_reg_ack_0 : boolean;
  signal addr_of_376_final_reg_req_1 : boolean;
  signal addr_of_376_final_reg_ack_1 : boolean;
  signal type_cast_718_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_660_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_660_inst_req_1 : boolean;
  signal type_cast_380_inst_req_0 : boolean;
  signal type_cast_380_inst_ack_0 : boolean;
  signal type_cast_380_inst_req_1 : boolean;
  signal type_cast_380_inst_ack_1 : boolean;
  signal type_cast_718_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_660_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_660_inst_req_0 : boolean;
  signal type_cast_646_inst_ack_1 : boolean;
  signal ptr_deref_383_store_0_req_0 : boolean;
  signal type_cast_646_inst_req_1 : boolean;
  signal ptr_deref_383_store_0_ack_0 : boolean;
  signal ptr_deref_383_store_0_req_1 : boolean;
  signal ptr_deref_383_store_0_ack_1 : boolean;
  signal type_cast_572_inst_ack_1 : boolean;
  signal type_cast_646_inst_ack_0 : boolean;
  signal type_cast_646_inst_req_0 : boolean;
  signal type_cast_572_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_642_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_642_inst_req_1 : boolean;
  signal ptr_deref_400_load_0_req_0 : boolean;
  signal ptr_deref_400_load_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_611_inst_ack_1 : boolean;
  signal ptr_deref_400_load_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_642_inst_ack_0 : boolean;
  signal ptr_deref_400_load_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_642_inst_req_0 : boolean;
  signal type_cast_572_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_req_0 : boolean;
  signal type_cast_700_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_ack_0 : boolean;
  signal type_cast_572_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_ack_1 : boolean;
  signal type_cast_736_inst_ack_1 : boolean;
  signal if_stmt_410_branch_req_0 : boolean;
  signal if_stmt_410_branch_ack_1 : boolean;
  signal if_stmt_410_branch_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_611_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_696_inst_ack_0 : boolean;
  signal type_cast_700_inst_req_1 : boolean;
  signal type_cast_736_inst_req_1 : boolean;
  signal STORE_pad_431_store_0_req_0 : boolean;
  signal STORE_pad_431_store_0_ack_0 : boolean;
  signal STORE_pad_431_store_0_req_1 : boolean;
  signal type_cast_628_inst_ack_1 : boolean;
  signal STORE_pad_431_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_435_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_435_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_435_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_435_inst_ack_1 : boolean;
  signal type_cast_439_inst_req_0 : boolean;
  signal type_cast_439_inst_ack_0 : boolean;
  signal type_cast_439_inst_req_1 : boolean;
  signal type_cast_439_inst_ack_1 : boolean;
  signal ptr_deref_450_store_0_req_0 : boolean;
  signal ptr_deref_450_store_0_ack_0 : boolean;
  signal ptr_deref_450_store_0_req_1 : boolean;
  signal ptr_deref_450_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_454_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_454_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_454_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_454_inst_ack_1 : boolean;
  signal type_cast_458_inst_req_0 : boolean;
  signal type_cast_458_inst_ack_0 : boolean;
  signal type_cast_458_inst_req_1 : boolean;
  signal type_cast_458_inst_ack_1 : boolean;
  signal ptr_deref_469_store_0_req_0 : boolean;
  signal ptr_deref_469_store_0_ack_0 : boolean;
  signal ptr_deref_469_store_0_req_1 : boolean;
  signal ptr_deref_469_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_473_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_473_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_473_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_473_inst_ack_1 : boolean;
  signal type_cast_477_inst_req_0 : boolean;
  signal type_cast_477_inst_ack_0 : boolean;
  signal type_cast_477_inst_req_1 : boolean;
  signal type_cast_477_inst_ack_1 : boolean;
  signal ptr_deref_488_store_0_req_0 : boolean;
  signal ptr_deref_488_store_0_ack_0 : boolean;
  signal ptr_deref_488_store_0_req_1 : boolean;
  signal ptr_deref_488_store_0_ack_1 : boolean;
  signal ptr_deref_501_load_0_req_0 : boolean;
  signal ptr_deref_501_load_0_ack_0 : boolean;
  signal ptr_deref_501_load_0_req_1 : boolean;
  signal ptr_deref_501_load_0_ack_1 : boolean;
  signal ptr_deref_513_load_0_req_0 : boolean;
  signal ptr_deref_513_load_0_ack_0 : boolean;
  signal ptr_deref_513_load_0_req_1 : boolean;
  signal ptr_deref_513_load_0_ack_1 : boolean;
  signal if_stmt_758_branch_req_0 : boolean;
  signal if_stmt_758_branch_ack_1 : boolean;
  signal if_stmt_758_branch_ack_0 : boolean;
  signal type_cast_769_inst_req_0 : boolean;
  signal type_cast_769_inst_ack_0 : boolean;
  signal type_cast_769_inst_req_1 : boolean;
  signal type_cast_769_inst_ack_1 : boolean;
  signal type_cast_350_inst_req_0 : boolean;
  signal type_cast_350_inst_ack_0 : boolean;
  signal type_cast_350_inst_req_1 : boolean;
  signal type_cast_350_inst_ack_1 : boolean;
  signal phi_stmt_347_req_0 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal phi_stmt_354_req_0 : boolean;
  signal phi_stmt_347_req_1 : boolean;
  signal type_cast_359_inst_req_0 : boolean;
  signal type_cast_359_inst_ack_0 : boolean;
  signal type_cast_359_inst_req_1 : boolean;
  signal type_cast_359_inst_ack_1 : boolean;
  signal phi_stmt_354_req_1 : boolean;
  signal phi_stmt_347_ack_0 : boolean;
  signal phi_stmt_354_ack_0 : boolean;
  signal type_cast_420_inst_req_0 : boolean;
  signal type_cast_420_inst_ack_0 : boolean;
  signal type_cast_420_inst_req_1 : boolean;
  signal type_cast_420_inst_ack_1 : boolean;
  signal phi_stmt_417_req_0 : boolean;
  signal phi_stmt_417_ack_0 : boolean;
  signal type_cast_427_inst_req_0 : boolean;
  signal type_cast_427_inst_ack_0 : boolean;
  signal type_cast_427_inst_req_1 : boolean;
  signal type_cast_427_inst_ack_1 : boolean;
  signal phi_stmt_424_req_0 : boolean;
  signal type_cast_429_inst_req_0 : boolean;
  signal type_cast_429_inst_ack_0 : boolean;
  signal type_cast_429_inst_req_1 : boolean;
  signal type_cast_429_inst_ack_1 : boolean;
  signal phi_stmt_424_req_1 : boolean;
  signal phi_stmt_424_ack_0 : boolean;
  signal phi_stmt_595_req_0 : boolean;
  signal type_cast_601_inst_req_0 : boolean;
  signal type_cast_601_inst_ack_0 : boolean;
  signal type_cast_601_inst_req_1 : boolean;
  signal type_cast_601_inst_ack_1 : boolean;
  signal phi_stmt_595_req_1 : boolean;
  signal phi_stmt_595_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_684_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_684: Block -- control-path 
    signal testConfigure_CP_684_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    testConfigure_CP_684_elements(0) <= testConfigure_CP_684_start;
    testConfigure_CP_684_symbol <= testConfigure_CP_684_elements(126);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	14 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/branch_block_stmt_283__entry__
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_update_start_
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_update_start_
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/ptr_deref_291_Split/split_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/ptr_deref_291_Split/split_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_update_start_
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337__entry__
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_update_start_
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/ptr_deref_291_Split/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/ptr_deref_291_Split/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_update_start_
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_root_address_calculated
      -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => RPIPE_zeropad_input_pipe_296_inst_req_0); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_300_inst_req_1); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_291_store_0_req_1); -- 
    cr_887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_317_inst_req_1); -- 
    rr_770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_291_store_0_req_0); -- 
    cr_859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_309_store_0_req_1); -- 
    cr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_326_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	19 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Sample/word_access_start/$exit
      -- 
    ra_771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_291_store_0_ack_0, ack => testConfigure_CP_684_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	21 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_Update/$exit
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_291_store_0_ack_1, ack => testConfigure_CP_684_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_update_start_
      -- CP-element group 3: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Update/$entry
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_296_inst_ack_0, ack => testConfigure_CP_684_elements(3)); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(3), ack => RPIPE_zeropad_input_pipe_296_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_296_Update/$exit
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_296_inst_ack_1, ack => testConfigure_CP_684_elements(4)); -- 
    rr_868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(4), ack => RPIPE_zeropad_input_pipe_313_inst_req_0); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(4), ack => type_cast_300_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_sample_completed_
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_300_inst_ack_0, ack => testConfigure_CP_684_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_300_update_completed_
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_300_inst_ack_1, ack => testConfigure_CP_684_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/ptr_deref_309_Split/split_req
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/ptr_deref_309_Split/$exit
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/ptr_deref_309_Split/$entry
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/word_access_start/word_0/rr
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/ptr_deref_309_Split/split_ack
      -- 
    rr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(7), ack => ptr_deref_309_store_0_req_0); -- 
    testConfigure_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(19) & testConfigure_CP_684_elements(6);
      gj_testConfigure_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	20 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Sample/word_access_start/$exit
      -- 
    ra_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_store_0_ack_0, ack => testConfigure_CP_684_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	21 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_Update/$exit
      -- 
    ca_860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_store_0_ack_1, ack => testConfigure_CP_684_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_update_start_
      -- CP-element group 10: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Update/cr
      -- 
    ra_869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_313_inst_ack_0, ack => testConfigure_CP_684_elements(10)); -- 
    cr_873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(10), ack => RPIPE_zeropad_input_pipe_313_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_313_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Sample/$entry
      -- 
    ca_874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_313_inst_ack_1, ack => testConfigure_CP_684_elements(11)); -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(11), ack => RPIPE_zeropad_input_pipe_336_inst_req_0); -- 
    rr_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(11), ack => type_cast_317_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Sample/ra
      -- 
    ra_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_0, ack => testConfigure_CP_684_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/type_cast_317_update_completed_
      -- 
    ca_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_1, ack => testConfigure_CP_684_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	0 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/ptr_deref_326_Split/$entry
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/ptr_deref_326_Split/$exit
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/word_access_start/word_0/rr
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/ptr_deref_326_Split/split_ack
      -- CP-element group 14: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/ptr_deref_326_Split/split_req
      -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(14), ack => ptr_deref_326_store_0_req_0); -- 
    testConfigure_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(20) & testConfigure_CP_684_elements(13);
      gj_testConfigure_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_sample_completed_
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_326_store_0_ack_0, ack => testConfigure_CP_684_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_326_Update/word_access_complete/word_0/$exit
      -- 
    ca_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_326_store_0_ack_1, ack => testConfigure_CP_684_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_update_start_
      -- CP-element group 17: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Update/cr
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_336_inst_ack_0, ack => testConfigure_CP_684_elements(17)); -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(17), ack => RPIPE_zeropad_input_pipe_336_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/RPIPE_zeropad_input_pipe_336_Update/ca
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_336_inst_ack_1, ack => testConfigure_CP_684_elements(18)); -- 
    -- CP-element group 19:  transition  delay-element  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	1 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	7 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_291_ptr_deref_309_delay
      -- 
    -- Element group testConfigure_CP_684_elements(19) is a control-delay.
    cp_element_19_delay: control_delay_element  generic map(name => " 19_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(1), ack => testConfigure_CP_684_elements(19), clk => clk, reset =>reset);
    -- CP-element group 20:  transition  delay-element  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	8 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/ptr_deref_309_ptr_deref_326_delay
      -- 
    -- Element group testConfigure_CP_684_elements(20) is a control-delay.
    cp_element_20_delay: control_delay_element  generic map(name => " 20_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(8), ack => testConfigure_CP_684_elements(20), clk => clk, reset =>reset);
    -- CP-element group 21:  branch  join  transition  place  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	9 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (10) 
      -- CP-element group 21: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337/$exit
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338__entry__
      -- CP-element group 21: 	 branch_block_stmt_283/assign_stmt_289_to_assign_stmt_337__exit__
      -- CP-element group 21: 	 branch_block_stmt_283/R_cmp87_339_place
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338_eval_test/$exit
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338_eval_test/branch_req
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338_dead_link/$entry
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338_else_link/$entry
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338_eval_test/$entry
      -- CP-element group 21: 	 branch_block_stmt_283/if_stmt_338_if_link/$entry
      -- 
    branch_req_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(21), ack => if_stmt_338_branch_req_0); -- 
    testConfigure_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(18) & testConfigure_CP_684_elements(9) & testConfigure_CP_684_elements(16) & testConfigure_CP_684_elements(2);
      gj_testConfigure_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  place  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	147 
    -- CP-element group 22: 	148 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_283/if_stmt_338_if_link/$exit
      -- CP-element group 22: 	 branch_block_stmt_283/if_stmt_338_if_link/if_choice_transition
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Update/cr
      -- 
    if_choice_transition_967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_338_branch_ack_1, ack => testConfigure_CP_684_elements(22)); -- 
    rr_2170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(22), ack => type_cast_427_inst_req_0); -- 
    cr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(22), ack => type_cast_427_inst_req_1); -- 
    -- CP-element group 23:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	134 
    -- CP-element group 23: 	135 
    -- CP-element group 23: 	136 
    -- CP-element group 23:  members (22) 
      -- CP-element group 23: 	 branch_block_stmt_283/entry_forx_xbodyx_xpreheader
      -- CP-element group 23: 	 branch_block_stmt_283/if_stmt_338_else_link/else_choice_transition
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 23: 	 branch_block_stmt_283/merge_stmt_344__exit__
      -- CP-element group 23: 	 branch_block_stmt_283/if_stmt_338_else_link/$exit
      -- CP-element group 23: 	 branch_block_stmt_283/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_283/merge_stmt_344_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_283/merge_stmt_344_PhiAck/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/merge_stmt_344_PhiAck/$exit
      -- CP-element group 23: 	 branch_block_stmt_283/merge_stmt_344_PhiAck/dummy
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_347/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Update/cr
      -- 
    else_choice_transition_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_338_branch_ack_0, ack => testConfigure_CP_684_elements(23)); -- 
    rr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(23), ack => type_cast_359_inst_req_0); -- 
    cr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(23), ack => type_cast_359_inst_req_1); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	142 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Sample/ra
      -- 
    ra_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_369_inst_ack_0, ack => testConfigure_CP_684_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	142 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	41 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Update/ca
      -- 
    ca_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_369_inst_ack_1, ack => testConfigure_CP_684_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	142 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	41 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_sample_complete
      -- CP-element group 26: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Sample/ack
      -- 
    ack_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_375_index_offset_ack_0, ack => testConfigure_CP_684_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	142 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (11) 
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_root_address_calculated
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_offset_calculated
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Update/ack
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_base_plus_offset/$entry
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_base_plus_offset/$exit
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_base_plus_offset/sum_rename_req
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_base_plus_offset/sum_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_request/$entry
      -- CP-element group 27: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_request/req
      -- 
    ack_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_375_index_offset_ack_1, ack => testConfigure_CP_684_elements(27)); -- 
    req_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(27), ack => addr_of_376_final_reg_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_request/$exit
      -- CP-element group 28: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_request/ack
      -- 
    ack_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_376_final_reg_ack_0, ack => testConfigure_CP_684_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	142 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (19) 
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_complete/$exit
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_complete/ack
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_word_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_root_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_address_resized
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_addr_resize/$entry
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_addr_resize/$exit
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_addr_resize/base_resize_req
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_addr_resize/base_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_plus_offset/$entry
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_plus_offset/$exit
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_plus_offset/sum_rename_req
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_base_plus_offset/sum_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_word_addrgen/$entry
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_word_addrgen/$exit
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_word_addrgen/root_register_req
      -- CP-element group 29: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_word_addrgen/root_register_ack
      -- 
    ack_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_376_final_reg_ack_1, ack => testConfigure_CP_684_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	142 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Sample/ra
      -- 
    ra_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_0, ack => testConfigure_CP_684_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	142 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Update/ca
      -- 
    ca_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_1, ack => testConfigure_CP_684_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/ptr_deref_383_Split/$entry
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/ptr_deref_383_Split/$exit
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/ptr_deref_383_Split/split_req
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/ptr_deref_383_Split/split_ack
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/word_access_start/$entry
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/word_access_start/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/word_access_start/word_0/rr
      -- 
    rr_1088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(32), ack => ptr_deref_383_store_0_req_0); -- 
    testConfigure_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(29) & testConfigure_CP_684_elements(31);
      gj_testConfigure_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	40 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Sample/word_access_start/word_0/ra
      -- 
    ra_1089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_383_store_0_ack_0, ack => testConfigure_CP_684_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	142 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/word_access_complete/word_0/ca
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_383_store_0_ack_1, ack => testConfigure_CP_684_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	40 
    -- CP-element group 35: 	142 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/word_access_start/$entry
      -- CP-element group 35: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/word_access_start/word_0/rr
      -- 
    rr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(35), ack => ptr_deref_400_load_0_req_0); -- 
    testConfigure_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(40) & testConfigure_CP_684_elements(142);
      gj_testConfigure_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/word_access_start/$exit
      -- CP-element group 36: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/word_access_start/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Sample/word_access_start/word_0/ra
      -- 
    ra_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_400_load_0_ack_0, ack => testConfigure_CP_684_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	142 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	41 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/word_access_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/word_access_complete/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/word_access_complete/word_0/ca
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/ptr_deref_400_Merge/$entry
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/ptr_deref_400_Merge/$exit
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/ptr_deref_400_Merge/merge_req
      -- CP-element group 37: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/ptr_deref_400_Merge/merge_ack
      -- 
    ca_1145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_400_load_0_ack_1, ack => testConfigure_CP_684_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	142 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_update_start_
      -- CP-element group 38: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Update/cr
      -- 
    ra_1159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_408_inst_ack_0, ack => testConfigure_CP_684_elements(38)); -- 
    cr_1163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(38), ack => RPIPE_zeropad_input_pipe_408_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Update/ca
      -- 
    ca_1164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_408_inst_ack_1, ack => testConfigure_CP_684_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	33 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	35 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_ptr_deref_400_delay
      -- 
    -- Element group testConfigure_CP_684_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(33), ack => testConfigure_CP_684_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  branch  join  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	25 
    -- CP-element group 41: 	26 
    -- CP-element group 41: 	34 
    -- CP-element group 41: 	37 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (10) 
      -- CP-element group 41: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/$exit
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410__entry__
      -- CP-element group 41: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409__exit__
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410_dead_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410_eval_test/$entry
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410_eval_test/$exit
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410_eval_test/branch_req
      -- CP-element group 41: 	 branch_block_stmt_283/R_cmp_411_place
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410_if_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_283/if_stmt_410_else_link/$entry
      -- 
    branch_req_1173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(41), ack => if_stmt_410_branch_req_0); -- 
    testConfigure_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(25) & testConfigure_CP_684_elements(26) & testConfigure_CP_684_elements(34) & testConfigure_CP_684_elements(37) & testConfigure_CP_684_elements(39);
      gj_testConfigure_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  place  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	127 
    -- CP-element group 42: 	128 
    -- CP-element group 42: 	130 
    -- CP-element group 42: 	131 
    -- CP-element group 42:  members (20) 
      -- CP-element group 42: 	 branch_block_stmt_283/if_stmt_410_if_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_283/if_stmt_410_if_link/if_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Update/cr
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Update/cr
      -- 
    if_choice_transition_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_410_branch_ack_1, ack => testConfigure_CP_684_elements(42)); -- 
    rr_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(42), ack => type_cast_350_inst_req_0); -- 
    cr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(42), ack => type_cast_350_inst_req_1); -- 
    rr_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(42), ack => type_cast_357_inst_req_0); -- 
    cr_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(42), ack => type_cast_357_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  place  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	143 
    -- CP-element group 43: 	144 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_283/if_stmt_410_else_link/$exit
      -- CP-element group 43: 	 branch_block_stmt_283/if_stmt_410_else_link/else_choice_transition
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_410_branch_ack_0, ack => testConfigure_CP_684_elements(43)); -- 
    rr_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(43), ack => type_cast_420_inst_req_0); -- 
    cr_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(43), ack => type_cast_420_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	154 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/word_access_start/$exit
      -- CP-element group 44: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/word_access_start/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/word_access_start/word_0/ra
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_431_store_0_ack_0, ack => testConfigure_CP_684_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	154 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	78 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/word_access_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/word_access_complete/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/word_access_complete/word_0/ca
      -- 
    ca_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_431_store_0_ack_1, ack => testConfigure_CP_684_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	154 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_update_start_
      -- CP-element group 46: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Update/cr
      -- 
    ra_1229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_435_inst_ack_0, ack => testConfigure_CP_684_elements(46)); -- 
    cr_1233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(46), ack => RPIPE_zeropad_input_pipe_435_inst_req_1); -- 
    -- CP-element group 47:  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	53 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Sample/rr
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Sample/rr
      -- 
    ca_1234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_435_inst_ack_1, ack => testConfigure_CP_684_elements(47)); -- 
    rr_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(47), ack => type_cast_439_inst_req_0); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(47), ack => RPIPE_zeropad_input_pipe_454_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Sample/ra
      -- 
    ra_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_439_inst_ack_0, ack => testConfigure_CP_684_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	154 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Update/ca
      -- 
    ca_1248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_439_inst_ack_1, ack => testConfigure_CP_684_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	154 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/ptr_deref_450_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/ptr_deref_450_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/ptr_deref_450_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/ptr_deref_450_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/word_access_start/word_0/rr
      -- 
    rr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(50), ack => ptr_deref_450_store_0_req_0); -- 
    testConfigure_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(49) & testConfigure_CP_684_elements(154);
      gj_testConfigure_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	76 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Sample/word_access_start/word_0/ra
      -- 
    ra_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_450_store_0_ack_0, ack => testConfigure_CP_684_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	154 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	78 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/word_access_complete/word_0/ca
      -- 
    ca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_450_store_0_ack_1, ack => testConfigure_CP_684_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	47 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_update_start_
      -- CP-element group 53: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Update/cr
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_454_inst_ack_0, ack => testConfigure_CP_684_elements(53)); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(53), ack => RPIPE_zeropad_input_pipe_454_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	60 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_454_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Sample/rr
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_454_inst_ack_1, ack => testConfigure_CP_684_elements(54)); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(54), ack => type_cast_458_inst_req_0); -- 
    rr_1384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(54), ack => RPIPE_zeropad_input_pipe_473_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Sample/ra
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_0, ack => testConfigure_CP_684_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	154 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Update/ca
      -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_1, ack => testConfigure_CP_684_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: 	76 
    -- CP-element group 57: 	154 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/ptr_deref_469_Split/$entry
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/ptr_deref_469_Split/$exit
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/ptr_deref_469_Split/split_req
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/ptr_deref_469_Split/split_ack
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/word_access_start/$entry
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/word_access_start/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/word_access_start/word_0/rr
      -- 
    rr_1364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(57), ack => ptr_deref_469_store_0_req_0); -- 
    testConfigure_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(56) & testConfigure_CP_684_elements(76) & testConfigure_CP_684_elements(154);
      gj_testConfigure_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	77 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/word_access_start/$exit
      -- CP-element group 58: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/word_access_start/word_0/$exit
      -- CP-element group 58: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Sample/word_access_start/word_0/ra
      -- 
    ra_1365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_469_store_0_ack_0, ack => testConfigure_CP_684_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	154 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	78 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/word_access_complete/$exit
      -- CP-element group 59: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/word_access_complete/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/word_access_complete/word_0/ca
      -- 
    ca_1376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_469_store_0_ack_1, ack => testConfigure_CP_684_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	54 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_update_start_
      -- CP-element group 60: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Sample/ra
      -- CP-element group 60: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Update/cr
      -- 
    ra_1385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_473_inst_ack_0, ack => testConfigure_CP_684_elements(60)); -- 
    cr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(60), ack => RPIPE_zeropad_input_pipe_473_inst_req_1); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_473_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Sample/rr
      -- 
    ca_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_473_inst_ack_1, ack => testConfigure_CP_684_elements(61)); -- 
    rr_1398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(61), ack => type_cast_477_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Sample/ra
      -- 
    ra_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_477_inst_ack_0, ack => testConfigure_CP_684_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	154 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Update/ca
      -- 
    ca_1404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_477_inst_ack_1, ack => testConfigure_CP_684_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: 	77 
    -- CP-element group 64: 	154 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/ptr_deref_488_Split/$entry
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/ptr_deref_488_Split/$exit
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/ptr_deref_488_Split/split_req
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/ptr_deref_488_Split/split_ack
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/word_access_start/word_0/rr
      -- 
    rr_1442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(64), ack => ptr_deref_488_store_0_req_0); -- 
    testConfigure_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(63) & testConfigure_CP_684_elements(77) & testConfigure_CP_684_elements(154);
      gj_testConfigure_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Sample/word_access_start/word_0/ra
      -- 
    ra_1443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_488_store_0_ack_0, ack => testConfigure_CP_684_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	154 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	78 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/word_access_complete/word_0/ca
      -- 
    ca_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_488_store_0_ack_1, ack => testConfigure_CP_684_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	154 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (5) 
      -- CP-element group 67: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/word_access_start/$exit
      -- CP-element group 67: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/word_access_start/word_0/$exit
      -- CP-element group 67: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/word_access_start/word_0/ra
      -- 
    ra_1488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_0_ack_0, ack => testConfigure_CP_684_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	154 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	73 
    -- CP-element group 68:  members (9) 
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/word_access_complete/$exit
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/word_access_complete/word_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/word_access_complete/word_0/ca
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/ptr_deref_501_Merge/$entry
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/ptr_deref_501_Merge/$exit
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/ptr_deref_501_Merge/merge_req
      -- CP-element group 68: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/ptr_deref_501_Merge/merge_ack
      -- 
    ca_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_0_ack_1, ack => testConfigure_CP_684_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	154 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/word_access_start/$exit
      -- CP-element group 69: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/word_access_start/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/word_access_start/word_0/ra
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_0_ack_0, ack => testConfigure_CP_684_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	154 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (9) 
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/word_access_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/word_access_complete/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/word_access_complete/word_0/ca
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/ptr_deref_513_Merge/$entry
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/ptr_deref_513_Merge/$exit
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/ptr_deref_513_Merge/merge_req
      -- CP-element group 70: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/ptr_deref_513_Merge/merge_ack
      -- 
    ca_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_0_ack_1, ack => testConfigure_CP_684_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	154 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/word_access_start/word_0/ra
      -- CP-element group 71: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/word_access_start/word_0/$exit
      -- CP-element group 71: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/word_access_start/$exit
      -- CP-element group 71: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_sample_completed_
      -- 
    ra_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_525_load_0_ack_0, ack => testConfigure_CP_684_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	154 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (9) 
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/ptr_deref_525_Merge/$exit
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/word_access_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/word_access_complete/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/word_access_complete/word_0/ca
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/ptr_deref_525_Merge/$entry
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/ptr_deref_525_Merge/merge_req
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/ptr_deref_525_Merge/merge_ack
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_update_completed_
      -- 
    ca_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_525_load_0_ack_1, ack => testConfigure_CP_684_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	68 
    -- CP-element group 73: 	70 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Sample/$entry
      -- 
    rr_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(73), ack => type_cast_539_inst_req_0); -- 
    testConfigure_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(68) & testConfigure_CP_684_elements(70) & testConfigure_CP_684_elements(72);
      gj_testConfigure_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_sample_completed_
      -- 
    ra_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_0, ack => testConfigure_CP_684_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	154 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_update_completed_
      -- 
    ca_1618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_1, ack => testConfigure_CP_684_elements(75)); -- 
    -- CP-element group 76:  transition  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	51 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	57 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_ptr_deref_469_delay
      -- 
    -- Element group testConfigure_CP_684_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(51), ack => testConfigure_CP_684_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	58 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	64 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_ptr_deref_488_delay
      -- 
    -- Element group testConfigure_CP_684_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(58), ack => testConfigure_CP_684_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  branch  join  transition  place  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	45 
    -- CP-element group 78: 	52 
    -- CP-element group 78: 	59 
    -- CP-element group 78: 	66 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (10) 
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553_eval_test/$entry
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553__entry__
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553_if_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553_eval_test/$exit
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553_eval_test/branch_req
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553_else_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552__exit__
      -- CP-element group 78: 	 branch_block_stmt_283/if_stmt_553_dead_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_283/R_cmp2684_554_place
      -- CP-element group 78: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/$exit
      -- 
    branch_req_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(78), ack => if_stmt_553_branch_req_0); -- 
    testConfigure_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(45) & testConfigure_CP_684_elements(52) & testConfigure_CP_684_elements(59) & testConfigure_CP_684_elements(66) & testConfigure_CP_684_elements(75);
      gj_testConfigure_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  place  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	161 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_283/if_stmt_553_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_283/if_stmt_553_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_283/forx_xend_forx_xend79
      -- CP-element group 79: 	 branch_block_stmt_283/forx_xend_forx_xend79_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_283/forx_xend_forx_xend79_PhiReq/$exit
      -- 
    if_choice_transition_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_553_branch_ack_1, ack => testConfigure_CP_684_elements(79)); -- 
    -- CP-element group 80:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (18) 
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_update_start_
      -- CP-element group 80: 	 branch_block_stmt_283/if_stmt_553_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/$entry
      -- CP-element group 80: 	 branch_block_stmt_283/if_stmt_553_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592__entry__
      -- CP-element group 80: 	 branch_block_stmt_283/merge_stmt_559__exit__
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_283/forx_xend_bbx_xnph
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_283/forx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_283/forx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_283/merge_stmt_559_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_283/merge_stmt_559_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_283/merge_stmt_559_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_283/merge_stmt_559_PhiAck/dummy
      -- 
    else_choice_transition_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_553_branch_ack_0, ack => testConfigure_CP_684_elements(80)); -- 
    cr_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(80), ack => type_cast_572_inst_req_1); -- 
    rr_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(80), ack => type_cast_572_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Sample/$exit
      -- 
    ra_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_572_inst_ack_0, ack => testConfigure_CP_684_elements(81)); -- 
    -- CP-element group 82:  transition  place  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	155 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28
      -- CP-element group 82: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592__exit__
      -- CP-element group 82: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/$exit
      -- CP-element group 82: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_283/assign_stmt_564_to_assign_stmt_592/type_cast_572_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/$entry
      -- CP-element group 82: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/phi_stmt_595/$entry
      -- CP-element group 82: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/$entry
      -- 
    ca_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_572_inst_ack_1, ack => testConfigure_CP_684_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	160 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	122 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Sample/ack
      -- CP-element group 83: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_sample_complete
      -- 
    ack_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_607_index_offset_ack_0, ack => testConfigure_CP_684_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	160 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (11) 
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Update/ack
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_base_plus_offset/$entry
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_base_plus_offset/$exit
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_base_plus_offset/sum_rename_req
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_base_plus_offset/sum_rename_ack
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_request/$entry
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_request/req
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_offset_calculated
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_root_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_sample_start_
      -- 
    ack_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_607_index_offset_ack_1, ack => testConfigure_CP_684_elements(84)); -- 
    req_1699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(84), ack => addr_of_608_final_reg_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_request/$exit
      -- CP-element group 85: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_request/ack
      -- CP-element group 85: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_sample_completed_
      -- 
    ack_1700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_608_final_reg_ack_0, ack => testConfigure_CP_684_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	160 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	119 
    -- CP-element group 86:  members (19) 
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_word_addrgen/$entry
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_word_addrgen/$exit
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_addr_resize/base_resize_req
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_address_calculated
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_complete/$exit
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_plus_offset/$entry
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_plus_offset/$exit
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_complete/ack
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_addr_resize/base_resize_ack
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_addr_resize/$exit
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_word_addrgen/root_register_ack
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_plus_offset/sum_rename_req
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_word_addrgen/root_register_req
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_plus_offset/sum_rename_ack
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_addr_resize/$entry
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_base_address_resized
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_root_address_calculated
      -- CP-element group 86: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_word_address_calculated
      -- 
    ack_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_608_final_reg_ack_1, ack => testConfigure_CP_684_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	160 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_update_start_
      -- CP-element group 87: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Update/$entry
      -- 
    ra_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_611_inst_ack_0, ack => testConfigure_CP_684_elements(87)); -- 
    cr_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(87), ack => RPIPE_zeropad_input_pipe_611_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	91 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Update/$exit
      -- 
    ca_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_611_inst_ack_1, ack => testConfigure_CP_684_elements(88)); -- 
    rr_1727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(88), ack => type_cast_615_inst_req_0); -- 
    rr_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(88), ack => RPIPE_zeropad_input_pipe_624_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_sample_completed_
      -- 
    ra_1728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_0, ack => testConfigure_CP_684_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	160 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	119 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_update_completed_
      -- 
    ca_1733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_1, ack => testConfigure_CP_684_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_update_start_
      -- CP-element group 91: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Update/cr
      -- 
    ra_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_624_inst_ack_0, ack => testConfigure_CP_684_elements(91)); -- 
    cr_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(91), ack => RPIPE_zeropad_input_pipe_624_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_624_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_sample_start_
      -- 
    ca_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_624_inst_ack_1, ack => testConfigure_CP_684_elements(92)); -- 
    rr_1755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(92), ack => type_cast_628_inst_req_0); -- 
    rr_1769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(92), ack => RPIPE_zeropad_input_pipe_642_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Sample/ra
      -- 
    ra_1756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_628_inst_ack_0, ack => testConfigure_CP_684_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	160 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	119 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Update/ca
      -- 
    ca_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_628_inst_ack_1, ack => testConfigure_CP_684_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Update/cr
      -- CP-element group 95: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_update_start_
      -- CP-element group 95: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_sample_completed_
      -- 
    ra_1770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_642_inst_ack_0, ack => testConfigure_CP_684_elements(95)); -- 
    cr_1774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(95), ack => RPIPE_zeropad_input_pipe_642_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_642_update_completed_
      -- 
    ca_1775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_642_inst_ack_1, ack => testConfigure_CP_684_elements(96)); -- 
    rr_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(96), ack => type_cast_646_inst_req_0); -- 
    rr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(96), ack => RPIPE_zeropad_input_pipe_660_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_sample_completed_
      -- 
    ra_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_646_inst_ack_0, ack => testConfigure_CP_684_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	160 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	119 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Update/ca
      -- CP-element group 98: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_update_completed_
      -- 
    ca_1789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_646_inst_ack_1, ack => testConfigure_CP_684_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Update/cr
      -- CP-element group 99: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_update_start_
      -- CP-element group 99: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_sample_completed_
      -- 
    ra_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_660_inst_ack_0, ack => testConfigure_CP_684_elements(99)); -- 
    cr_1802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(99), ack => RPIPE_zeropad_input_pipe_660_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_660_update_completed_
      -- 
    ca_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_660_inst_ack_1, ack => testConfigure_CP_684_elements(100)); -- 
    rr_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(100), ack => type_cast_664_inst_req_0); -- 
    rr_1825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(100), ack => RPIPE_zeropad_input_pipe_678_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_sample_completed_
      -- 
    ra_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_0, ack => testConfigure_CP_684_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	160 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	119 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_update_completed_
      -- 
    ca_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_1, ack => testConfigure_CP_684_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_update_start_
      -- CP-element group 103: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_sample_completed_
      -- 
    ra_1826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_678_inst_ack_0, ack => testConfigure_CP_684_elements(103)); -- 
    cr_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(103), ack => RPIPE_zeropad_input_pipe_678_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_678_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Sample/$entry
      -- 
    ca_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_678_inst_ack_1, ack => testConfigure_CP_684_elements(104)); -- 
    rr_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(104), ack => type_cast_682_inst_req_0); -- 
    rr_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(104), ack => RPIPE_zeropad_input_pipe_696_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Sample/ra
      -- 
    ra_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_682_inst_ack_0, ack => testConfigure_CP_684_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	160 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	119 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Update/ca
      -- 
    ca_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_682_inst_ack_1, ack => testConfigure_CP_684_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_update_start_
      -- CP-element group 107: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Sample/ra
      -- 
    ra_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_696_inst_ack_0, ack => testConfigure_CP_684_elements(107)); -- 
    cr_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(107), ack => RPIPE_zeropad_input_pipe_696_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_696_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_sample_start_
      -- 
    ca_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_696_inst_ack_1, ack => testConfigure_CP_684_elements(108)); -- 
    rr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(108), ack => type_cast_700_inst_req_0); -- 
    rr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(108), ack => RPIPE_zeropad_input_pipe_714_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Sample/$exit
      -- 
    ra_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_700_inst_ack_0, ack => testConfigure_CP_684_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	160 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	119 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Update/$exit
      -- 
    ca_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_700_inst_ack_1, ack => testConfigure_CP_684_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_update_start_
      -- CP-element group 111: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_sample_completed_
      -- 
    ra_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_714_inst_ack_0, ack => testConfigure_CP_684_elements(111)); -- 
    cr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(111), ack => RPIPE_zeropad_input_pipe_714_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_714_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Sample/$entry
      -- 
    ca_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_714_inst_ack_1, ack => testConfigure_CP_684_elements(112)); -- 
    rr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(112), ack => type_cast_718_inst_req_0); -- 
    rr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(112), ack => RPIPE_zeropad_input_pipe_732_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Sample/$exit
      -- 
    ra_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_718_inst_ack_0, ack => testConfigure_CP_684_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	160 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	119 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Update/$exit
      -- 
    ca_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_718_inst_ack_1, ack => testConfigure_CP_684_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_update_start_
      -- CP-element group 115: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Update/$entry
      -- 
    ra_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_732_inst_ack_0, ack => testConfigure_CP_684_elements(115)); -- 
    cr_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => RPIPE_zeropad_input_pipe_732_inst_req_1); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_732_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_sample_start_
      -- 
    ca_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_732_inst_ack_1, ack => testConfigure_CP_684_elements(116)); -- 
    rr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(116), ack => type_cast_736_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_sample_completed_
      -- 
    ra_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_736_inst_ack_0, ack => testConfigure_CP_684_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	160 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Update/ca
      -- 
    ca_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_736_inst_ack_1, ack => testConfigure_CP_684_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	86 
    -- CP-element group 119: 	90 
    -- CP-element group 119: 	94 
    -- CP-element group 119: 	98 
    -- CP-element group 119: 	102 
    -- CP-element group 119: 	106 
    -- CP-element group 119: 	110 
    -- CP-element group 119: 	114 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (9) 
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/ptr_deref_744_Split/$entry
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/ptr_deref_744_Split/$exit
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/ptr_deref_744_Split/split_ack
      -- CP-element group 119: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/ptr_deref_744_Split/split_req
      -- 
    rr_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(119), ack => ptr_deref_744_store_0_req_0); -- 
    testConfigure_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(86) & testConfigure_CP_684_elements(90) & testConfigure_CP_684_elements(94) & testConfigure_CP_684_elements(98) & testConfigure_CP_684_elements(102) & testConfigure_CP_684_elements(106) & testConfigure_CP_684_elements(110) & testConfigure_CP_684_elements(114) & testConfigure_CP_684_elements(118);
      gj_testConfigure_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/word_access_start/word_0/ra
      -- CP-element group 120: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Sample/word_access_start/$exit
      -- 
    ra_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_744_store_0_ack_0, ack => testConfigure_CP_684_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	160 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/word_access_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/word_access_complete/word_0/$exit
      -- 
    ca_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_744_store_0_ack_1, ack => testConfigure_CP_684_elements(121)); -- 
    -- CP-element group 122:  branch  join  transition  place  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	83 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (10) 
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758__entry__
      -- CP-element group 122: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757__exit__
      -- CP-element group 122: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/$exit
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758_dead_link/$entry
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758_eval_test/$entry
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758_eval_test/$exit
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758_eval_test/branch_req
      -- CP-element group 122: 	 branch_block_stmt_283/R_exitcond10_759_place
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758_if_link/$entry
      -- CP-element group 122: 	 branch_block_stmt_283/if_stmt_758_else_link/$entry
      -- 
    branch_req_1987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(122), ack => if_stmt_758_branch_req_0); -- 
    testConfigure_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(83) & testConfigure_CP_684_elements(121);
      gj_testConfigure_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  transition  place  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	161 
    -- CP-element group 123:  members (13) 
      -- CP-element group 123: 	 branch_block_stmt_283/forx_xend79x_xloopexit_forx_xend79
      -- CP-element group 123: 	 branch_block_stmt_283/merge_stmt_764__exit__
      -- CP-element group 123: 	 branch_block_stmt_283/if_stmt_758_if_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_283/if_stmt_758_if_link/if_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_283/forx_xbody28_forx_xend79x_xloopexit
      -- CP-element group 123: 	 branch_block_stmt_283/forx_xbody28_forx_xend79x_xloopexit_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_283/forx_xbody28_forx_xend79x_xloopexit_PhiReq/$exit
      -- CP-element group 123: 	 branch_block_stmt_283/merge_stmt_764_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_283/merge_stmt_764_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_283/merge_stmt_764_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_283/merge_stmt_764_PhiAck/dummy
      -- CP-element group 123: 	 branch_block_stmt_283/forx_xend79x_xloopexit_forx_xend79_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_283/forx_xend79x_xloopexit_forx_xend79_PhiReq/$exit
      -- 
    if_choice_transition_1992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_758_branch_ack_1, ack => testConfigure_CP_684_elements(123)); -- 
    -- CP-element group 124:  fork  transition  place  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	156 
    -- CP-element group 124: 	157 
    -- CP-element group 124:  members (12) 
      -- CP-element group 124: 	 branch_block_stmt_283/if_stmt_758_else_link/$exit
      -- CP-element group 124: 	 branch_block_stmt_283/if_stmt_758_else_link/else_choice_transition
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Sample/rr
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_758_branch_ack_0, ack => testConfigure_CP_684_elements(124)); -- 
    rr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(124), ack => type_cast_601_inst_req_0); -- 
    cr_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(124), ack => type_cast_601_inst_req_1); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	161 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Sample/ra
      -- 
    ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_0, ack => testConfigure_CP_684_elements(125)); -- 
    -- CP-element group 126:  transition  place  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	161 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (16) 
      -- CP-element group 126: 	 branch_block_stmt_283/$exit
      -- CP-element group 126: 	 $exit
      -- CP-element group 126: 	 branch_block_stmt_283/return__
      -- CP-element group 126: 	 branch_block_stmt_283/assign_stmt_770__exit__
      -- CP-element group 126: 	 branch_block_stmt_283/merge_stmt_772__exit__
      -- CP-element group 126: 	 branch_block_stmt_283/branch_block_stmt_283__exit__
      -- CP-element group 126: 	 branch_block_stmt_283/assign_stmt_770/$exit
      -- CP-element group 126: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Update/ca
      -- CP-element group 126: 	 branch_block_stmt_283/return___PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_283/return___PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_283/merge_stmt_772_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_283/merge_stmt_772_PhiAck/$entry
      -- CP-element group 126: 	 branch_block_stmt_283/merge_stmt_772_PhiAck/$exit
      -- CP-element group 126: 	 branch_block_stmt_283/merge_stmt_772_PhiAck/dummy
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_1, ack => testConfigure_CP_684_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	42 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Sample/ra
      -- 
    ra_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_350_inst_ack_0, ack => testConfigure_CP_684_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	42 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/Update/ca
      -- 
    ca_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_350_inst_ack_1, ack => testConfigure_CP_684_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/$exit
      -- CP-element group 129: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/$exit
      -- CP-element group 129: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/$exit
      -- CP-element group 129: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_350/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_req
      -- 
    phi_stmt_347_req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_347_req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(129), ack => phi_stmt_347_req_0); -- 
    testConfigure_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(127) & testConfigure_CP_684_elements(128);
      gj_testConfigure_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	42 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Sample/ra
      -- 
    ra_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => testConfigure_CP_684_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	42 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/Update/ca
      -- 
    ca_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => testConfigure_CP_684_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/$exit
      -- CP-element group 132: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/$exit
      -- CP-element group 132: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/$exit
      -- CP-element group 132: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_357/SplitProtocol/$exit
      -- CP-element group 132: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_req
      -- 
    phi_stmt_354_req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_354_req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(132), ack => phi_stmt_354_req_0); -- 
    testConfigure_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(130) & testConfigure_CP_684_elements(131);
      gj_testConfigure_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	129 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	139 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_283/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(129) & testConfigure_CP_684_elements(132);
      gj_testConfigure_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  output  delay-element  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	23 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	138 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_347/$exit
      -- CP-element group 134: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/$exit
      -- CP-element group 134: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_sources/type_cast_353_konst_delay_trans
      -- CP-element group 134: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_347/phi_stmt_347_req
      -- 
    phi_stmt_347_req_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_347_req_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(134), ack => phi_stmt_347_req_1); -- 
    -- Element group testConfigure_CP_684_elements(134) is a control-delay.
    cp_element_134_delay: control_delay_element  generic map(name => " 134_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(23), ack => testConfigure_CP_684_elements(134), clk => clk, reset =>reset);
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	23 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Sample/ra
      -- 
    ra_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_0, ack => testConfigure_CP_684_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	23 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/Update/ca
      -- 
    ca_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_1, ack => testConfigure_CP_684_elements(136)); -- 
    -- CP-element group 137:  join  transition  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (5) 
      -- CP-element group 137: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/$exit
      -- CP-element group 137: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/$exit
      -- CP-element group 137: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/$exit
      -- CP-element group 137: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_sources/type_cast_359/SplitProtocol/$exit
      -- CP-element group 137: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_354/phi_stmt_354_req
      -- 
    phi_stmt_354_req_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_354_req_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(137), ack => phi_stmt_354_req_1); -- 
    testConfigure_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(135) & testConfigure_CP_684_elements(136);
      gj_testConfigure_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	134 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_283/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(134) & testConfigure_CP_684_elements(137);
      gj_testConfigure_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  merge  fork  transition  place  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	133 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_283/merge_stmt_346_PhiReqMerge
      -- CP-element group 139: 	 branch_block_stmt_283/merge_stmt_346_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(139) <= OrReduce(testConfigure_CP_684_elements(133) & testConfigure_CP_684_elements(138));
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_283/merge_stmt_346_PhiAck/phi_stmt_347_ack
      -- 
    phi_stmt_347_ack_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_347_ack_0, ack => testConfigure_CP_684_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_283/merge_stmt_346_PhiAck/phi_stmt_354_ack
      -- 
    phi_stmt_354_ack_2116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_354_ack_0, ack => testConfigure_CP_684_elements(141)); -- 
    -- CP-element group 142:  join  fork  transition  place  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	24 
    -- CP-element group 142: 	25 
    -- CP-element group 142: 	26 
    -- CP-element group 142: 	27 
    -- CP-element group 142: 	29 
    -- CP-element group 142: 	30 
    -- CP-element group 142: 	31 
    -- CP-element group 142: 	34 
    -- CP-element group 142: 	35 
    -- CP-element group 142: 	37 
    -- CP-element group 142: 	38 
    -- CP-element group 142:  members (64) 
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_update_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_369_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409__entry__
      -- CP-element group 142: 	 branch_block_stmt_283/merge_stmt_346__exit__
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_update_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_resized_1
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_scaled_1
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_computed_1
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_resize_1/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_resize_1/$exit
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_resize_1/index_resize_req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_resize_1/index_resize_ack
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_scale_1/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_scale_1/$exit
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_scale_1/scale_rename_req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_index_scale_1/scale_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_update_start
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Sample/req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/array_obj_ref_375_final_index_sum_regn_Update/req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_complete/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/addr_of_376_complete/req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_update_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/type_cast_380_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_update_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/word_access_complete/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/word_access_complete/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_383_Update/word_access_complete/word_0/cr
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_update_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_word_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_root_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_address_resized
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_addr_resize/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_addr_resize/$exit
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_addr_resize/base_resize_req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_addr_resize/base_resize_ack
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_plus_offset/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_plus_offset/$exit
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_plus_offset/sum_rename_req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_base_plus_offset/sum_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_word_addrgen/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_word_addrgen/$exit
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_word_addrgen/root_register_req
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_word_addrgen/root_register_ack
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/word_access_complete/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/word_access_complete/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/ptr_deref_400_Update/word_access_complete/word_0/cr
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_283/assign_stmt_366_to_assign_stmt_409/RPIPE_zeropad_input_pipe_408_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_283/merge_stmt_346_PhiAck/$exit
      -- 
    rr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => type_cast_369_inst_req_0); -- 
    cr_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => type_cast_369_inst_req_1); -- 
    req_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => array_obj_ref_375_index_offset_req_0); -- 
    req_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => array_obj_ref_375_index_offset_req_1); -- 
    req_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => addr_of_376_final_reg_req_1); -- 
    rr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => type_cast_380_inst_req_0); -- 
    cr_1049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => type_cast_380_inst_req_1); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => ptr_deref_383_store_0_req_1); -- 
    cr_1144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => ptr_deref_400_load_0_req_1); -- 
    rr_1158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(142), ack => RPIPE_zeropad_input_pipe_408_inst_req_0); -- 
    testConfigure_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(140) & testConfigure_CP_684_elements(141);
      gj_testConfigure_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	43 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Sample/ra
      -- 
    ra_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_420_inst_ack_0, ack => testConfigure_CP_684_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	43 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/Update/ca
      -- 
    ca_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_420_inst_ack_1, ack => testConfigure_CP_684_elements(144)); -- 
    -- CP-element group 145:  join  transition  place  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (8) 
      -- CP-element group 145: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 145: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/$exit
      -- CP-element group 145: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/$exit
      -- CP-element group 145: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/$exit
      -- CP-element group 145: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_sources/type_cast_420/SplitProtocol/$exit
      -- CP-element group 145: 	 branch_block_stmt_283/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_417/phi_stmt_417_req
      -- CP-element group 145: 	 branch_block_stmt_283/merge_stmt_416_PhiReqMerge
      -- CP-element group 145: 	 branch_block_stmt_283/merge_stmt_416_PhiAck/$entry
      -- 
    phi_stmt_417_req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_417_req_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(145), ack => phi_stmt_417_req_0); -- 
    testConfigure_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(143) & testConfigure_CP_684_elements(144);
      gj_testConfigure_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	150 
    -- CP-element group 146: 	151 
    -- CP-element group 146:  members (13) 
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend
      -- CP-element group 146: 	 branch_block_stmt_283/merge_stmt_416__exit__
      -- CP-element group 146: 	 branch_block_stmt_283/merge_stmt_416_PhiAck/$exit
      -- CP-element group 146: 	 branch_block_stmt_283/merge_stmt_416_PhiAck/phi_stmt_417_ack
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Update/cr
      -- 
    phi_stmt_417_ack_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_417_ack_0, ack => testConfigure_CP_684_elements(146)); -- 
    rr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(146), ack => type_cast_429_inst_req_0); -- 
    cr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(146), ack => type_cast_429_inst_req_1); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	22 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Sample/ra
      -- 
    ra_2171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_427_inst_ack_0, ack => testConfigure_CP_684_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	22 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/Update/ca
      -- 
    ca_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_427_inst_ack_1, ack => testConfigure_CP_684_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	153 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/$exit
      -- CP-element group 149: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/$exit
      -- CP-element group 149: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/$exit
      -- CP-element group 149: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/$exit
      -- CP-element group 149: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_427/SplitProtocol/$exit
      -- CP-element group 149: 	 branch_block_stmt_283/entry_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_req
      -- 
    phi_stmt_424_req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_424_req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(149), ack => phi_stmt_424_req_0); -- 
    testConfigure_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(147) & testConfigure_CP_684_elements(148);
      gj_testConfigure_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	146 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Sample/ra
      -- 
    ra_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_429_inst_ack_0, ack => testConfigure_CP_684_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	146 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/Update/ca
      -- 
    ca_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_429_inst_ack_1, ack => testConfigure_CP_684_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 152: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/$exit
      -- CP-element group 152: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/$exit
      -- CP-element group 152: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/$exit
      -- CP-element group 152: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_sources/type_cast_429/SplitProtocol/$exit
      -- CP-element group 152: 	 branch_block_stmt_283/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_424/phi_stmt_424_req
      -- 
    phi_stmt_424_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_424_req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(152), ack => phi_stmt_424_req_1); -- 
    testConfigure_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(150) & testConfigure_CP_684_elements(151);
      gj_testConfigure_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  merge  transition  place  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	149 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_283/merge_stmt_423_PhiReqMerge
      -- CP-element group 153: 	 branch_block_stmt_283/merge_stmt_423_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(153) <= OrReduce(testConfigure_CP_684_elements(149) & testConfigure_CP_684_elements(152));
    -- CP-element group 154:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	44 
    -- CP-element group 154: 	45 
    -- CP-element group 154: 	46 
    -- CP-element group 154: 	49 
    -- CP-element group 154: 	50 
    -- CP-element group 154: 	52 
    -- CP-element group 154: 	56 
    -- CP-element group 154: 	57 
    -- CP-element group 154: 	59 
    -- CP-element group 154: 	63 
    -- CP-element group 154: 	64 
    -- CP-element group 154: 	66 
    -- CP-element group 154: 	67 
    -- CP-element group 154: 	68 
    -- CP-element group 154: 	69 
    -- CP-element group 154: 	70 
    -- CP-element group 154: 	71 
    -- CP-element group 154: 	72 
    -- CP-element group 154: 	75 
    -- CP-element group 154:  members (177) 
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/word_access_start/word_0/rr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552__entry__
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/word_access_start/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/merge_stmt_423__exit__
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Sample/word_access_start/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_word_addrgen/root_register_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_539_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/STORE_pad_431_Split/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/STORE_pad_431_Split/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/STORE_pad_431_Split/split_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/STORE_pad_431_Split/split_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/word_access_start/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/word_access_start/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Sample/word_access_start/word_0/rr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/STORE_pad_431_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/RPIPE_zeropad_input_pipe_435_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_439_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_word_addrgen/root_register_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_450_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_458_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_word_addrgen/root_register_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_469_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/type_cast_477_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_word_addrgen/root_register_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_488_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_word_addrgen/root_register_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/word_access_start/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/word_access_start/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Sample/word_access_start/word_0/rr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_501_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_word_addrgen/root_register_ack
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/word_access_start/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/word_access_start/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Sample/word_access_start/word_0/rr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/word_access_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/word_access_complete/word_0/$entry
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_513_Update/word_access_complete/word_0/cr
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_update_start_
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_283/assign_stmt_433_to_assign_stmt_552/ptr_deref_525_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_283/merge_stmt_423_PhiAck/$exit
      -- CP-element group 154: 	 branch_block_stmt_283/merge_stmt_423_PhiAck/phi_stmt_424_ack
      -- 
    phi_stmt_424_ack_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_424_ack_0, ack => testConfigure_CP_684_elements(154)); -- 
    cr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_525_load_0_req_1); -- 
    rr_1587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_525_load_0_req_0); -- 
    cr_1617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => type_cast_539_inst_req_1); -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => STORE_pad_431_store_0_req_0); -- 
    cr_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => STORE_pad_431_store_0_req_1); -- 
    rr_1228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => RPIPE_zeropad_input_pipe_435_inst_req_0); -- 
    cr_1247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => type_cast_439_inst_req_1); -- 
    cr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_450_store_0_req_1); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => type_cast_458_inst_req_1); -- 
    cr_1375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_469_store_0_req_1); -- 
    cr_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => type_cast_477_inst_req_1); -- 
    cr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_488_store_0_req_1); -- 
    rr_1487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_501_load_0_req_0); -- 
    cr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_501_load_0_req_1); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_513_load_0_req_0); -- 
    cr_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(154), ack => ptr_deref_513_load_0_req_1); -- 
    -- CP-element group 155:  transition  output  delay-element  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	82 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	159 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/$exit
      -- CP-element group 155: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/phi_stmt_595/$exit
      -- CP-element group 155: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/$exit
      -- CP-element group 155: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_599_konst_delay_trans
      -- CP-element group 155: 	 branch_block_stmt_283/bbx_xnph_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_req
      -- 
    phi_stmt_595_req_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_595_req_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(155), ack => phi_stmt_595_req_0); -- 
    -- Element group testConfigure_CP_684_elements(155) is a control-delay.
    cp_element_155_delay: control_delay_element  generic map(name => " 155_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(82), ack => testConfigure_CP_684_elements(155), clk => clk, reset =>reset);
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	124 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Sample/ra
      -- 
    ra_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_0, ack => testConfigure_CP_684_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	124 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (2) 
      -- CP-element group 157: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/Update/ca
      -- 
    ca_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_1, ack => testConfigure_CP_684_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/$exit
      -- CP-element group 158: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/$exit
      -- CP-element group 158: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/$exit
      -- CP-element group 158: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/$exit
      -- CP-element group 158: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_sources/type_cast_601/SplitProtocol/$exit
      -- CP-element group 158: 	 branch_block_stmt_283/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_595/phi_stmt_595_req
      -- 
    phi_stmt_595_req_2257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_595_req_2257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(158), ack => phi_stmt_595_req_1); -- 
    testConfigure_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(156) & testConfigure_CP_684_elements(157);
      gj_testConfigure_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  merge  transition  place  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	155 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_283/merge_stmt_594_PhiReqMerge
      -- CP-element group 159: 	 branch_block_stmt_283/merge_stmt_594_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(159) <= OrReduce(testConfigure_CP_684_elements(155) & testConfigure_CP_684_elements(158));
    -- CP-element group 160:  fork  transition  place  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	83 
    -- CP-element group 160: 	84 
    -- CP-element group 160: 	86 
    -- CP-element group 160: 	87 
    -- CP-element group 160: 	90 
    -- CP-element group 160: 	94 
    -- CP-element group 160: 	98 
    -- CP-element group 160: 	102 
    -- CP-element group 160: 	106 
    -- CP-element group 160: 	110 
    -- CP-element group 160: 	114 
    -- CP-element group 160: 	118 
    -- CP-element group 160: 	121 
    -- CP-element group 160:  members (56) 
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/word_access_complete/word_0/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Update/req
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Sample/rr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_update_start
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_scale_1/scale_rename_ack
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_computed_1
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_682_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_resize_1/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Sample/req
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757__entry__
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_scale_1/$exit
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_scale_1/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_resize_1/index_resize_req
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_complete/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_scale_1/scale_rename_req
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_final_index_sum_regn_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/merge_stmt_594__exit__
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_complete/req
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_resize_1/index_resize_ack
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_resize_1/$exit
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/RPIPE_zeropad_input_pipe_611_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/word_access_complete/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_628_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_664_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_scaled_1
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/array_obj_ref_607_index_resized_1
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/addr_of_608_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_718_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_615_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_646_update_start_
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/ptr_deref_744_Update/word_access_complete/word_0/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_736_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_283/assign_stmt_609_to_assign_stmt_757/type_cast_700_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_283/merge_stmt_594_PhiAck/$exit
      -- CP-element group 160: 	 branch_block_stmt_283/merge_stmt_594_PhiAck/phi_stmt_595_ack
      -- 
    phi_stmt_595_ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_595_ack_0, ack => testConfigure_CP_684_elements(160)); -- 
    cr_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => ptr_deref_744_store_0_req_1); -- 
    req_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => array_obj_ref_607_index_offset_req_1); -- 
    rr_1713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => RPIPE_zeropad_input_pipe_611_inst_req_0); -- 
    cr_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_682_inst_req_1); -- 
    cr_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_628_inst_req_1); -- 
    cr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_664_inst_req_1); -- 
    req_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => array_obj_ref_607_index_offset_req_0); -- 
    cr_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_615_inst_req_1); -- 
    req_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => addr_of_608_final_reg_req_1); -- 
    cr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_718_inst_req_1); -- 
    cr_1788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_646_inst_req_1); -- 
    cr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_700_inst_req_1); -- 
    cr_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(160), ack => type_cast_736_inst_req_1); -- 
    -- CP-element group 161:  merge  fork  transition  place  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	79 
    -- CP-element group 161: 	123 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	125 
    -- CP-element group 161: 	126 
    -- CP-element group 161:  members (13) 
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770__entry__
      -- CP-element group 161: 	 branch_block_stmt_283/merge_stmt_766__exit__
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/$entry
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_update_start_
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_283/assign_stmt_770/type_cast_769_Update/cr
      -- CP-element group 161: 	 branch_block_stmt_283/merge_stmt_766_PhiReqMerge
      -- CP-element group 161: 	 branch_block_stmt_283/merge_stmt_766_PhiAck/$entry
      -- CP-element group 161: 	 branch_block_stmt_283/merge_stmt_766_PhiAck/$exit
      -- CP-element group 161: 	 branch_block_stmt_283/merge_stmt_766_PhiAck/dummy
      -- 
    rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(161), ack => type_cast_769_inst_req_0); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(161), ack => type_cast_769_inst_req_1); -- 
    testConfigure_CP_684_elements(161) <= OrReduce(testConfigure_CP_684_elements(79) & testConfigure_CP_684_elements(123));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar97_374_resized : std_logic_vector(6 downto 0);
    signal R_indvar97_374_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_606_resized : std_logic_vector(13 downto 0);
    signal R_indvar_606_scaled : std_logic_vector(13 downto 0);
    signal STORE_pad_431_data_0 : std_logic_vector(7 downto 0);
    signal STORE_pad_431_word_address_0 : std_logic_vector(0 downto 0);
    signal add41_652 : std_logic_vector(63 downto 0);
    signal add47_670 : std_logic_vector(63 downto 0);
    signal add53_688 : std_logic_vector(63 downto 0);
    signal add59_706 : std_logic_vector(63 downto 0);
    signal add65_724 : std_logic_vector(63 downto 0);
    signal add71_742 : std_logic_vector(63 downto 0);
    signal add_634 : std_logic_vector(63 downto 0);
    signal array_obj_ref_375_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_375_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_375_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_375_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_375_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_375_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_607_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_607_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_607_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_607_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_607_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_607_root_address : std_logic_vector(13 downto 0);
    signal arrayidx75_609 : std_logic_vector(31 downto 0);
    signal arrayidx_377 : std_logic_vector(31 downto 0);
    signal call10_436 : std_logic_vector(7 downto 0);
    signal call12_455 : std_logic_vector(7 downto 0);
    signal call14_474 : std_logic_vector(7 downto 0);
    signal call1_314 : std_logic_vector(7 downto 0);
    signal call30_612 : std_logic_vector(7 downto 0);
    signal call33_625 : std_logic_vector(7 downto 0);
    signal call38_643 : std_logic_vector(7 downto 0);
    signal call44_661 : std_logic_vector(7 downto 0);
    signal call50_679 : std_logic_vector(7 downto 0);
    signal call56_697 : std_logic_vector(7 downto 0);
    signal call588_337 : std_logic_vector(7 downto 0);
    signal call590_354 : std_logic_vector(7 downto 0);
    signal call5_409 : std_logic_vector(7 downto 0);
    signal call5x_xlcssa1_417 : std_logic_vector(7 downto 0);
    signal call5x_xlcssa_424 : std_logic_vector(7 downto 0);
    signal call62_715 : std_logic_vector(7 downto 0);
    signal call68_733 : std_logic_vector(7 downto 0);
    signal call_297 : std_logic_vector(7 downto 0);
    signal cmp2684_552 : std_logic_vector(0 downto 0);
    signal cmp87_334 : std_logic_vector(0 downto 0);
    signal cmp_406 : std_logic_vector(0 downto 0);
    signal conv11_440 : std_logic_vector(31 downto 0);
    signal conv13_459 : std_logic_vector(31 downto 0);
    signal conv15_478 : std_logic_vector(31 downto 0);
    signal conv21_540 : std_logic_vector(63 downto 0);
    signal conv2_318 : std_logic_vector(31 downto 0);
    signal conv31_616 : std_logic_vector(63 downto 0);
    signal conv35_629 : std_logic_vector(63 downto 0);
    signal conv40_647 : std_logic_vector(63 downto 0);
    signal conv46_665 : std_logic_vector(63 downto 0);
    signal conv52_683 : std_logic_vector(63 downto 0);
    signal conv58_701 : std_logic_vector(63 downto 0);
    signal conv64_719 : std_logic_vector(63 downto 0);
    signal conv6_381 : std_logic_vector(31 downto 0);
    signal conv70_737 : std_logic_vector(63 downto 0);
    signal conv_301 : std_logic_vector(31 downto 0);
    signal exitcond10_757 : std_logic_vector(0 downto 0);
    signal iNsTr_0_289 : std_logic_vector(31 downto 0);
    signal iNsTr_12_448 : std_logic_vector(31 downto 0);
    signal iNsTr_15_467 : std_logic_vector(31 downto 0);
    signal iNsTr_18_486 : std_logic_vector(31 downto 0);
    signal iNsTr_20_498 : std_logic_vector(31 downto 0);
    signal iNsTr_21_510 : std_logic_vector(31 downto 0);
    signal iNsTr_22_522 : std_logic_vector(31 downto 0);
    signal iNsTr_28_397 : std_logic_vector(31 downto 0);
    signal iNsTr_3_307 : std_logic_vector(31 downto 0);
    signal iNsTr_6_324 : std_logic_vector(31 downto 0);
    signal inc_370 : std_logic_vector(31 downto 0);
    signal indvar97_347 : std_logic_vector(63 downto 0);
    signal indvar_595 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_752 : std_logic_vector(63 downto 0);
    signal mul20_536 : std_logic_vector(31 downto 0);
    signal mul_531 : std_logic_vector(31 downto 0);
    signal ptr_deref_291_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_291_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_291_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_291_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_291_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_291_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_309_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_309_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_309_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_309_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_309_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_309_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_326_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_326_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_326_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_326_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_326_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_326_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_383_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_383_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_383_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_383_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_383_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_383_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_400_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_400_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_400_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_400_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_400_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_450_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_450_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_450_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_450_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_450_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_450_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_469_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_469_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_469_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_469_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_469_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_469_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_488_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_488_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_488_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_488_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_488_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_488_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_501_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_501_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_501_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_501_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_501_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_513_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_513_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_513_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_513_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_513_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_525_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_525_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_525_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_525_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_525_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_744_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_744_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_744_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_744_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_744_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_744_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl37_640 : std_logic_vector(63 downto 0);
    signal shl43_658 : std_logic_vector(63 downto 0);
    signal shl49_676 : std_logic_vector(63 downto 0);
    signal shl55_694 : std_logic_vector(63 downto 0);
    signal shl61_712 : std_logic_vector(63 downto 0);
    signal shl67_730 : std_logic_vector(63 downto 0);
    signal shl_622 : std_logic_vector(63 downto 0);
    signal shr83x_xmask_546 : std_logic_vector(63 downto 0);
    signal tmp17_502 : std_logic_vector(31 downto 0);
    signal tmp18_514 : std_logic_vector(31 downto 0);
    signal tmp19_526 : std_logic_vector(31 downto 0);
    signal tmp3_401 : std_logic_vector(31 downto 0);
    signal tmp4_564 : std_logic_vector(31 downto 0);
    signal tmp5_569 : std_logic_vector(31 downto 0);
    signal tmp6_573 : std_logic_vector(63 downto 0);
    signal tmp7_579 : std_logic_vector(63 downto 0);
    signal tmp8_585 : std_logic_vector(0 downto 0);
    signal tmp99_391 : std_logic_vector(63 downto 0);
    signal tmp_366 : std_logic_vector(63 downto 0);
    signal type_cast_293_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_332_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_350_wire : std_logic_vector(63 downto 0);
    signal type_cast_353_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_357_wire : std_logic_vector(7 downto 0);
    signal type_cast_359_wire : std_logic_vector(7 downto 0);
    signal type_cast_364_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_389_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_420_wire : std_logic_vector(7 downto 0);
    signal type_cast_427_wire : std_logic_vector(7 downto 0);
    signal type_cast_429_wire : std_logic_vector(7 downto 0);
    signal type_cast_544_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_550_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_577_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_583_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_590_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_599_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_601_wire : std_logic_vector(63 downto 0);
    signal type_cast_620_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_638_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_656_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_674_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_692_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_710_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_728_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_750_wire_constant : std_logic_vector(63 downto 0);
    signal umax9_592 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_pad_431_word_address_0 <= "0";
    array_obj_ref_375_constant_part_of_offset <= "0000011";
    array_obj_ref_375_offset_scale_factor_0 <= "1000000";
    array_obj_ref_375_offset_scale_factor_1 <= "0000001";
    array_obj_ref_375_resized_base_address <= "0000000";
    array_obj_ref_607_constant_part_of_offset <= "00000000000000";
    array_obj_ref_607_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_607_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_607_resized_base_address <= "00000000000000";
    iNsTr_0_289 <= "00000000000000000000000000000000";
    iNsTr_12_448 <= "00000000000000000000000000000011";
    iNsTr_15_467 <= "00000000000000000000000000000100";
    iNsTr_18_486 <= "00000000000000000000000000000101";
    iNsTr_20_498 <= "00000000000000000000000000000011";
    iNsTr_21_510 <= "00000000000000000000000000000100";
    iNsTr_22_522 <= "00000000000000000000000000000101";
    iNsTr_28_397 <= "00000000000000000000000000000010";
    iNsTr_3_307 <= "00000000000000000000000000000001";
    iNsTr_6_324 <= "00000000000000000000000000000010";
    ptr_deref_291_word_offset_0 <= "0000000";
    ptr_deref_309_word_offset_0 <= "0000000";
    ptr_deref_326_word_offset_0 <= "0000000";
    ptr_deref_383_word_offset_0 <= "0000000";
    ptr_deref_400_word_offset_0 <= "0000000";
    ptr_deref_450_word_offset_0 <= "0000000";
    ptr_deref_469_word_offset_0 <= "0000000";
    ptr_deref_488_word_offset_0 <= "0000000";
    ptr_deref_501_word_offset_0 <= "0000000";
    ptr_deref_513_word_offset_0 <= "0000000";
    ptr_deref_525_word_offset_0 <= "0000000";
    ptr_deref_744_word_offset_0 <= "00000000000000";
    type_cast_293_wire_constant <= "00000000000000000000000000000101";
    type_cast_332_wire_constant <= "00000000";
    type_cast_353_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_389_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_544_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_550_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_577_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_583_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_590_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_599_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_620_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_638_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_656_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_674_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_692_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_710_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_728_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_750_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_347: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_350_wire & type_cast_353_wire_constant;
      req <= phi_stmt_347_req_0 & phi_stmt_347_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_347",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_347_ack_0,
          idata => idata,
          odata => indvar97_347,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_347
    phi_stmt_354: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_357_wire & type_cast_359_wire;
      req <= phi_stmt_354_req_0 & phi_stmt_354_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_354",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_354_ack_0,
          idata => idata,
          odata => call590_354,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_354
    phi_stmt_417: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_420_wire;
      req(0) <= phi_stmt_417_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_417",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_417_ack_0,
          idata => idata,
          odata => call5x_xlcssa1_417,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_417
    phi_stmt_424: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_427_wire & type_cast_429_wire;
      req <= phi_stmt_424_req_0 & phi_stmt_424_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_424",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_424_ack_0,
          idata => idata,
          odata => call5x_xlcssa_424,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_424
    phi_stmt_595: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_599_wire_constant & type_cast_601_wire;
      req <= phi_stmt_595_req_0 & phi_stmt_595_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_595",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_595_ack_0,
          idata => idata,
          odata => indvar_595,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_595
    -- flow-through select operator MUX_591_inst
    umax9_592 <= tmp7_579 when (tmp8_585(0) /=  '0') else type_cast_590_wire_constant;
    addr_of_376_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_376_final_reg_req_0;
      addr_of_376_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_376_final_reg_req_1;
      addr_of_376_final_reg_ack_1<= rack(0);
      addr_of_376_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_376_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_375_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_608_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_608_final_reg_req_0;
      addr_of_608_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_608_final_reg_req_1;
      addr_of_608_final_reg_ack_1<= rack(0);
      addr_of_608_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_608_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_607_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx75_609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_300_inst_req_0;
      type_cast_300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_300_inst_req_1;
      type_cast_300_inst_ack_1<= rack(0);
      type_cast_300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_317_inst_req_0;
      type_cast_317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_317_inst_req_1;
      type_cast_317_inst_ack_1<= rack(0);
      type_cast_317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_314,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_318,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_350_inst_req_0;
      type_cast_350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_350_inst_req_1;
      type_cast_350_inst_ack_1<= rack(0);
      type_cast_350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp99_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_350_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_357_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_359_inst_req_0;
      type_cast_359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_359_inst_req_1;
      type_cast_359_inst_ack_1<= rack(0);
      type_cast_359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call588_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_359_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_369_inst_req_0;
      type_cast_369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_369_inst_req_1;
      type_cast_369_inst_ack_1<= rack(0);
      type_cast_369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_369_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_380_inst_req_0;
      type_cast_380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_380_inst_req_1;
      type_cast_380_inst_ack_1<= rack(0);
      type_cast_380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call590_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_420_inst_req_0;
      type_cast_420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_420_inst_req_1;
      type_cast_420_inst_ack_1<= rack(0);
      type_cast_420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_420_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_427_inst_req_0;
      type_cast_427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_427_inst_req_1;
      type_cast_427_inst_ack_1<= rack(0);
      type_cast_427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call588_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_427_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_429_inst_req_0;
      type_cast_429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_429_inst_req_1;
      type_cast_429_inst_ack_1<= rack(0);
      type_cast_429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5x_xlcssa1_417,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_429_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_439_inst_req_0;
      type_cast_439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_439_inst_req_1;
      type_cast_439_inst_ack_1<= rack(0);
      type_cast_439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_440,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_458_inst_req_0;
      type_cast_458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_458_inst_req_1;
      type_cast_458_inst_ack_1<= rack(0);
      type_cast_458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call12_455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_459,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_477_inst_req_0;
      type_cast_477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_477_inst_req_1;
      type_cast_477_inst_ack_1<= rack(0);
      type_cast_477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_539_inst_req_0;
      type_cast_539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_539_inst_req_1;
      type_cast_539_inst_ack_1<= rack(0);
      type_cast_539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul20_536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_572_inst_req_0;
      type_cast_572_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_572_inst_req_1;
      type_cast_572_inst_ack_1<= rack(0);
      type_cast_572_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_572_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_573,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_601_inst_req_0;
      type_cast_601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_601_inst_req_1;
      type_cast_601_inst_ack_1<= rack(0);
      type_cast_601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_752,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_601_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_615_inst_req_0;
      type_cast_615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_615_inst_req_1;
      type_cast_615_inst_ack_1<= rack(0);
      type_cast_615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_628_inst_req_0;
      type_cast_628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_628_inst_req_1;
      type_cast_628_inst_ack_1<= rack(0);
      type_cast_628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_628_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call33_625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_629,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_646_inst_req_0;
      type_cast_646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_646_inst_req_1;
      type_cast_646_inst_ack_1<= rack(0);
      type_cast_646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_646_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call38_643,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_647,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_664_inst_req_0;
      type_cast_664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_664_inst_req_1;
      type_cast_664_inst_ack_1<= rack(0);
      type_cast_664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_682_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_682_inst_req_0;
      type_cast_682_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_682_inst_req_1;
      type_cast_682_inst_ack_1<= rack(0);
      type_cast_682_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_682_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_679,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_683,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_700_inst_req_0;
      type_cast_700_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_700_inst_req_1;
      type_cast_700_inst_ack_1<= rack(0);
      type_cast_700_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_700_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_697,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_701,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_718_inst_req_0;
      type_cast_718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_718_inst_req_1;
      type_cast_718_inst_ack_1<= rack(0);
      type_cast_718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_736_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_736_inst_req_0;
      type_cast_736_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_736_inst_req_1;
      type_cast_736_inst_ack_1<= rack(0);
      type_cast_736_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_736_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_737,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_769_inst_req_0;
      type_cast_769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_769_inst_req_1;
      type_cast_769_inst_ack_1<= rack(0);
      type_cast_769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul20_536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_pad_431_gather_scatter
    process(call5x_xlcssa_424) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call5x_xlcssa_424;
      ov(7 downto 0) := iv;
      STORE_pad_431_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_375_index_1_rename
    process(R_indvar97_374_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar97_374_resized;
      ov(6 downto 0) := iv;
      R_indvar97_374_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_375_index_1_resize
    process(indvar97_347) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar97_347;
      ov := iv(6 downto 0);
      R_indvar97_374_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_375_root_address_inst
    process(array_obj_ref_375_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_375_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_375_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_607_index_1_rename
    process(R_indvar_606_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_606_resized;
      ov(13 downto 0) := iv;
      R_indvar_606_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_607_index_1_resize
    process(indvar_595) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_595;
      ov := iv(13 downto 0);
      R_indvar_606_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_607_root_address_inst
    process(array_obj_ref_607_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_607_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_607_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_291_addr_0
    process(ptr_deref_291_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_291_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_291_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_291_base_resize
    process(iNsTr_0_289) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_289;
      ov := iv(6 downto 0);
      ptr_deref_291_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_291_gather_scatter
    process(type_cast_293_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_293_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_291_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_291_root_address_inst
    process(ptr_deref_291_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_291_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_291_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_309_addr_0
    process(ptr_deref_309_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_309_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_309_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_309_base_resize
    process(iNsTr_3_307) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_307;
      ov := iv(6 downto 0);
      ptr_deref_309_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_309_gather_scatter
    process(conv_301) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_301;
      ov(31 downto 0) := iv;
      ptr_deref_309_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_309_root_address_inst
    process(ptr_deref_309_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_309_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_309_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_326_addr_0
    process(ptr_deref_326_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_326_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_326_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_326_base_resize
    process(iNsTr_6_324) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_324;
      ov := iv(6 downto 0);
      ptr_deref_326_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_326_gather_scatter
    process(conv2_318) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv2_318;
      ov(31 downto 0) := iv;
      ptr_deref_326_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_326_root_address_inst
    process(ptr_deref_326_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_326_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_326_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_addr_0
    process(ptr_deref_383_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_383_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_base_resize
    process(arrayidx_377) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_377;
      ov := iv(6 downto 0);
      ptr_deref_383_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_gather_scatter
    process(conv6_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv6_381;
      ov(31 downto 0) := iv;
      ptr_deref_383_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_root_address_inst
    process(ptr_deref_383_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_383_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_400_addr_0
    process(ptr_deref_400_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_400_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_400_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_400_base_resize
    process(iNsTr_28_397) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_28_397;
      ov := iv(6 downto 0);
      ptr_deref_400_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_400_gather_scatter
    process(ptr_deref_400_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_400_data_0;
      ov(31 downto 0) := iv;
      tmp3_401 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_400_root_address_inst
    process(ptr_deref_400_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_400_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_400_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_450_addr_0
    process(ptr_deref_450_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_450_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_450_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_450_base_resize
    process(iNsTr_12_448) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_12_448;
      ov := iv(6 downto 0);
      ptr_deref_450_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_450_gather_scatter
    process(conv11_440) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv11_440;
      ov(31 downto 0) := iv;
      ptr_deref_450_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_450_root_address_inst
    process(ptr_deref_450_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_450_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_450_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_addr_0
    process(ptr_deref_469_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_469_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_469_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_base_resize
    process(iNsTr_15_467) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_467;
      ov := iv(6 downto 0);
      ptr_deref_469_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_gather_scatter
    process(conv13_459) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv13_459;
      ov(31 downto 0) := iv;
      ptr_deref_469_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_root_address_inst
    process(ptr_deref_469_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_469_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_469_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_addr_0
    process(ptr_deref_488_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_488_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_base_resize
    process(iNsTr_18_486) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_486;
      ov := iv(6 downto 0);
      ptr_deref_488_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_gather_scatter
    process(conv15_478) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv15_478;
      ov(31 downto 0) := iv;
      ptr_deref_488_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_root_address_inst
    process(ptr_deref_488_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_488_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_addr_0
    process(ptr_deref_501_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_501_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_501_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_base_resize
    process(iNsTr_20_498) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_20_498;
      ov := iv(6 downto 0);
      ptr_deref_501_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_gather_scatter
    process(ptr_deref_501_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_501_data_0;
      ov(31 downto 0) := iv;
      tmp17_502 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_root_address_inst
    process(ptr_deref_501_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_501_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_501_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_addr_0
    process(ptr_deref_513_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_513_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_513_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_base_resize
    process(iNsTr_21_510) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_510;
      ov := iv(6 downto 0);
      ptr_deref_513_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_gather_scatter
    process(ptr_deref_513_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_513_data_0;
      ov(31 downto 0) := iv;
      tmp18_514 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_root_address_inst
    process(ptr_deref_513_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_513_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_513_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_525_addr_0
    process(ptr_deref_525_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_525_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_525_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_525_base_resize
    process(iNsTr_22_522) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_22_522;
      ov := iv(6 downto 0);
      ptr_deref_525_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_525_gather_scatter
    process(ptr_deref_525_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_525_data_0;
      ov(31 downto 0) := iv;
      tmp19_526 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_525_root_address_inst
    process(ptr_deref_525_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_525_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_525_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_744_addr_0
    process(ptr_deref_744_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_744_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_744_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_744_base_resize
    process(arrayidx75_609) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx75_609;
      ov := iv(13 downto 0);
      ptr_deref_744_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_744_gather_scatter
    process(add71_742) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add71_742;
      ov(63 downto 0) := iv;
      ptr_deref_744_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_744_root_address_inst
    process(ptr_deref_744_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_744_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_744_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_338_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp87_334;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_338_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_338_branch_req_0,
          ack0 => if_stmt_338_branch_ack_0,
          ack1 => if_stmt_338_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_410_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_406;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_410_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_410_branch_req_0,
          ack0 => if_stmt_410_branch_ack_0,
          ack1 => if_stmt_410_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_553_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp2684_552;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_553_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_553_branch_req_0,
          ack0 => if_stmt_553_branch_ack_0,
          ack1 => if_stmt_553_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_758_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond10_757;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_758_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_758_branch_req_0,
          ack0 => if_stmt_758_branch_ack_0,
          ack1 => if_stmt_758_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_365_inst
    process(indvar97_347) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar97_347, type_cast_364_wire_constant, tmp_var);
      tmp_366 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_390_inst
    process(indvar97_347) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar97_347, type_cast_389_wire_constant, tmp_var);
      tmp99_391 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_751_inst
    process(indvar_595) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_595, type_cast_750_wire_constant, tmp_var);
      indvarx_xnext_752 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_545_inst
    process(conv21_540) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv21_540, type_cast_544_wire_constant, tmp_var);
      shr83x_xmask_546 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_551_inst
    process(shr83x_xmask_546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr83x_xmask_546, type_cast_550_wire_constant, tmp_var);
      cmp2684_552 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_756_inst
    process(indvarx_xnext_752, umax9_592) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_752, umax9_592, tmp_var);
      exitcond10_757 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_333_inst
    process(call1_314) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call1_314, type_cast_332_wire_constant, tmp_var);
      cmp87_334 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_578_inst
    process(tmp6_573) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp6_573, type_cast_577_wire_constant, tmp_var);
      tmp7_579 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_530_inst
    process(tmp18_514, tmp17_502) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp18_514, tmp17_502, tmp_var);
      mul_531 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_535_inst
    process(mul_531, tmp19_526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_531, tmp19_526, tmp_var);
      mul20_536 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_563_inst
    process(tmp18_514, tmp17_502) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp18_514, tmp17_502, tmp_var);
      tmp4_564 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_568_inst
    process(tmp4_564, tmp19_526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_564, tmp19_526, tmp_var);
      tmp5_569 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_633_inst
    process(shl_622, conv35_629) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_622, conv35_629, tmp_var);
      add_634 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_651_inst
    process(shl37_640, conv40_647) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl37_640, conv40_647, tmp_var);
      add41_652 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_669_inst
    process(shl43_658, conv46_665) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl43_658, conv46_665, tmp_var);
      add47_670 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_687_inst
    process(shl49_676, conv52_683) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl49_676, conv52_683, tmp_var);
      add53_688 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_705_inst
    process(shl55_694, conv58_701) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl55_694, conv58_701, tmp_var);
      add59_706 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_723_inst
    process(shl61_712, conv64_719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl61_712, conv64_719, tmp_var);
      add65_724 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_741_inst
    process(shl67_730, conv70_737) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl67_730, conv70_737, tmp_var);
      add71_742 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_621_inst
    process(conv31_616) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv31_616, type_cast_620_wire_constant, tmp_var);
      shl_622 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_639_inst
    process(add_634) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_634, type_cast_638_wire_constant, tmp_var);
      shl37_640 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_657_inst
    process(add41_652) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add41_652, type_cast_656_wire_constant, tmp_var);
      shl43_658 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_675_inst
    process(add47_670) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add47_670, type_cast_674_wire_constant, tmp_var);
      shl49_676 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_693_inst
    process(add53_688) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add53_688, type_cast_692_wire_constant, tmp_var);
      shl55_694 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_711_inst
    process(add59_706) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add59_706, type_cast_710_wire_constant, tmp_var);
      shl61_712 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_729_inst
    process(add65_724) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add65_724, type_cast_728_wire_constant, tmp_var);
      shl67_730 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_584_inst
    process(tmp7_579) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp7_579, type_cast_583_wire_constant, tmp_var);
      tmp8_585 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_405_inst
    process(inc_370, tmp3_401) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_370, tmp3_401, tmp_var);
      cmp_406 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_375_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar97_374_scaled;
      array_obj_ref_375_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_375_index_offset_req_0;
      array_obj_ref_375_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_375_index_offset_req_1;
      array_obj_ref_375_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_607_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_606_scaled;
      array_obj_ref_607_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_607_index_offset_req_0;
      array_obj_ref_607_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_607_index_offset_req_1;
      array_obj_ref_607_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_513_load_0 ptr_deref_525_load_0 ptr_deref_501_load_0 ptr_deref_400_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_513_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_525_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_501_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_400_load_0_req_0;
      ptr_deref_513_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_525_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_501_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_400_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_513_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_525_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_501_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_400_load_0_req_1;
      ptr_deref_513_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_525_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_501_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_400_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_513_word_address_0 & ptr_deref_525_word_address_0 & ptr_deref_501_word_address_0 & ptr_deref_400_word_address_0;
      ptr_deref_513_data_0 <= data_out(127 downto 96);
      ptr_deref_525_data_0 <= data_out(95 downto 64);
      ptr_deref_501_data_0 <= data_out(63 downto 32);
      ptr_deref_400_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_pad_431_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_pad_431_store_0_req_0;
      STORE_pad_431_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_pad_431_store_0_req_1;
      STORE_pad_431_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_pad_431_word_address_0;
      data_in <= STORE_pad_431_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(0 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_291_store_0 ptr_deref_309_store_0 ptr_deref_326_store_0 ptr_deref_383_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_291_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_309_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_326_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_383_store_0_req_0;
      ptr_deref_291_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_309_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_326_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_383_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_291_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_309_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_326_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_383_store_0_req_1;
      ptr_deref_291_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_309_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_326_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_383_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_291_word_address_0 & ptr_deref_309_word_address_0 & ptr_deref_326_word_address_0 & ptr_deref_383_word_address_0;
      data_in <= ptr_deref_291_data_0 & ptr_deref_309_data_0 & ptr_deref_326_data_0 & ptr_deref_383_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_450_store_0 ptr_deref_469_store_0 ptr_deref_488_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_450_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_469_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_488_store_0_req_0;
      ptr_deref_450_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_469_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_488_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_450_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_469_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_488_store_0_req_1;
      ptr_deref_450_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_469_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_488_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_450_word_address_0 & ptr_deref_469_word_address_0 & ptr_deref_488_word_address_0;
      data_in <= ptr_deref_450_data_0 & ptr_deref_469_data_0 & ptr_deref_488_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(6 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_744_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_744_store_0_req_0;
      ptr_deref_744_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_744_store_0_req_1;
      ptr_deref_744_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_744_word_address_0;
      data_in <= ptr_deref_744_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_696_inst RPIPE_zeropad_input_pipe_732_inst RPIPE_zeropad_input_pipe_714_inst RPIPE_zeropad_input_pipe_660_inst RPIPE_zeropad_input_pipe_611_inst RPIPE_zeropad_input_pipe_624_inst RPIPE_zeropad_input_pipe_678_inst RPIPE_zeropad_input_pipe_642_inst RPIPE_zeropad_input_pipe_296_inst RPIPE_zeropad_input_pipe_313_inst RPIPE_zeropad_input_pipe_336_inst RPIPE_zeropad_input_pipe_408_inst RPIPE_zeropad_input_pipe_435_inst RPIPE_zeropad_input_pipe_454_inst RPIPE_zeropad_input_pipe_473_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(119 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 14 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 14 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 14 downto 0);
      signal guard_vector : std_logic_vector( 14 downto 0);
      constant outBUFs : IntegerArray(14 downto 0) := (14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(14 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false);
      constant guardBuffering: IntegerArray(14 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2);
      -- 
    begin -- 
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_696_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_732_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_714_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_660_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_611_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_624_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_678_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_642_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_296_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_313_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_336_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_408_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_435_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_454_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_473_inst_req_0;
      RPIPE_zeropad_input_pipe_696_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_732_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_714_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_660_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_611_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_624_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_678_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_642_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_296_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_313_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_336_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_408_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_435_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_454_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_473_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_696_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_732_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_714_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_660_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_611_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_624_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_678_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_642_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_296_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_313_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_336_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_408_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_435_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_454_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_473_inst_req_1;
      RPIPE_zeropad_input_pipe_696_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_732_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_714_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_660_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_611_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_624_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_678_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_642_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_296_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_313_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_336_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_408_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_435_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_454_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_473_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      call56_697 <= data_out(119 downto 112);
      call68_733 <= data_out(111 downto 104);
      call62_715 <= data_out(103 downto 96);
      call44_661 <= data_out(95 downto 88);
      call30_612 <= data_out(87 downto 80);
      call33_625 <= data_out(79 downto 72);
      call50_679 <= data_out(71 downto 64);
      call38_643 <= data_out(63 downto 56);
      call_297 <= data_out(55 downto 48);
      call1_314 <= data_out(47 downto 40);
      call588_337 <= data_out(39 downto 32);
      call5_409 <= data_out(31 downto 24);
      call10_436 <= data_out(23 downto 16);
      call12_455 <= data_out(15 downto 8);
      call14_474 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 15, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 15,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_2294_start: Boolean;
  signal timer_CP_2294_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_778_load_0_req_0 : boolean;
  signal LOAD_count_778_load_0_ack_0 : boolean;
  signal LOAD_count_778_load_0_req_1 : boolean;
  signal LOAD_count_778_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_2294_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_2294_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_2294_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_2294_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_2294: Block -- control-path 
    signal timer_CP_2294_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_2294_elements(0) <= timer_CP_2294_start;
    timer_CP_2294_symbol <= timer_CP_2294_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_779/$entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Update/$entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_sample_start_
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_update_start_
      -- CP-element group 0: 	 assign_stmt_779/LOAD_count_778_Sample/word_access_start/word_0/$entry
      -- 
    rr_2315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_2294_elements(0), ack => LOAD_count_778_load_0_req_0); -- 
    cr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_2294_elements(0), ack => LOAD_count_778_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_779/LOAD_count_778_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_779/LOAD_count_778_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_779/LOAD_count_778_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_779/LOAD_count_778_sample_completed_
      -- CP-element group 1: 	 assign_stmt_779/LOAD_count_778_Sample/word_access_start/$exit
      -- 
    ra_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_778_load_0_ack_0, ack => timer_CP_2294_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_779/$exit
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/$exit
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_update_completed_
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/LOAD_count_778_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/LOAD_count_778_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/LOAD_count_778_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_779/LOAD_count_778_Update/LOAD_count_778_Merge/merge_ack
      -- 
    ca_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_778_load_0_ack_1, ack => timer_CP_2294_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_778_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_778_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_778_word_address_0 <= "0";
    -- equivalence LOAD_count_778_gather_scatter
    process(LOAD_count_778_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_778_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_778_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_778_load_0_req_0;
      LOAD_count_778_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_778_load_0_req_1;
      LOAD_count_778_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_778_word_address_0;
      LOAD_count_778_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    Block2_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_2450_start: Boolean;
  signal zeropad3D_CP_2450_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_803_call_req_0 : boolean;
  signal call_stmt_803_call_ack_0 : boolean;
  signal call_stmt_803_call_req_1 : boolean;
  signal call_stmt_803_call_ack_1 : boolean;
  signal call_stmt_806_call_req_0 : boolean;
  signal call_stmt_806_call_ack_0 : boolean;
  signal call_stmt_806_call_req_1 : boolean;
  signal call_stmt_806_call_ack_1 : boolean;
  signal type_cast_811_inst_req_0 : boolean;
  signal type_cast_811_inst_ack_0 : boolean;
  signal type_cast_811_inst_req_1 : boolean;
  signal type_cast_811_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_813_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_813_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_813_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_813_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_816_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_816_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_816_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_816_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_819_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_819_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_819_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_819_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_822_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_822_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_822_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_822_inst_ack_1 : boolean;
  signal RPIPE_Block0_complete_826_inst_req_0 : boolean;
  signal RPIPE_Block0_complete_826_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_826_inst_req_1 : boolean;
  signal RPIPE_Block0_complete_826_inst_ack_1 : boolean;
  signal RPIPE_Block1_complete_829_inst_req_0 : boolean;
  signal RPIPE_Block1_complete_829_inst_ack_0 : boolean;
  signal RPIPE_Block1_complete_829_inst_req_1 : boolean;
  signal RPIPE_Block1_complete_829_inst_ack_1 : boolean;
  signal RPIPE_Block2_complete_832_inst_req_0 : boolean;
  signal RPIPE_Block2_complete_832_inst_ack_0 : boolean;
  signal RPIPE_Block2_complete_832_inst_req_1 : boolean;
  signal RPIPE_Block2_complete_832_inst_ack_1 : boolean;
  signal RPIPE_Block3_complete_835_inst_req_0 : boolean;
  signal RPIPE_Block3_complete_835_inst_ack_0 : boolean;
  signal RPIPE_Block3_complete_835_inst_req_1 : boolean;
  signal RPIPE_Block3_complete_835_inst_ack_1 : boolean;
  signal call_stmt_839_call_req_0 : boolean;
  signal call_stmt_839_call_ack_0 : boolean;
  signal call_stmt_839_call_req_1 : boolean;
  signal call_stmt_839_call_ack_1 : boolean;
  signal type_cast_843_inst_req_0 : boolean;
  signal type_cast_843_inst_ack_0 : boolean;
  signal type_cast_843_inst_req_1 : boolean;
  signal type_cast_843_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_850_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_850_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_850_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_850_inst_ack_1 : boolean;
  signal call_stmt_854_call_req_0 : boolean;
  signal call_stmt_854_call_ack_0 : boolean;
  signal call_stmt_854_call_req_1 : boolean;
  signal call_stmt_854_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_2450_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2450_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_2450_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2450_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_2450: Block -- control-path 
    signal zeropad3D_CP_2450_elements: BooleanArray(31 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_2450_elements(0) <= zeropad3D_CP_2450_start;
    zeropad3D_CP_2450_symbol <= zeropad3D_CP_2450_elements(31);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_801/$entry
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/$entry
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_update_start_
      -- CP-element group 0: 	 branch_block_stmt_801/branch_block_stmt_801__entry__
      -- CP-element group 0: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Update/$entry
      -- 
    crr_2478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(0), ack => call_stmt_803_call_req_0); -- 
    ccr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(0), ack => call_stmt_803_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_sample_completed_
      -- 
    cra_2479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_803_call_ack_0, ack => zeropad3D_CP_2450_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (40) 
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_803/$exit
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_update_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_update_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_803__exit__
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Update/ccr
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836__entry__
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_803/call_stmt_803_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Sample/rr
      -- 
    cca_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_803_call_ack_1, ack => zeropad3D_CP_2450_elements(2)); -- 
    crr_2495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => call_stmt_806_call_req_0); -- 
    ccr_2500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => call_stmt_806_call_req_1); -- 
    cr_2514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => type_cast_811_inst_req_1); -- 
    req_2523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => WPIPE_Block0_starting_813_inst_req_0); -- 
    req_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => WPIPE_Block1_starting_816_inst_req_0); -- 
    req_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => WPIPE_Block2_starting_819_inst_req_0); -- 
    req_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => WPIPE_Block3_starting_822_inst_req_0); -- 
    rr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => RPIPE_Block0_complete_826_inst_req_0); -- 
    rr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => RPIPE_Block1_complete_829_inst_req_0); -- 
    rr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => RPIPE_Block2_complete_832_inst_req_0); -- 
    rr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(2), ack => RPIPE_Block3_complete_835_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Sample/$exit
      -- 
    cra_2496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_806_call_ack_0, ack => zeropad3D_CP_2450_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/call_stmt_806_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Sample/rr
      -- 
    cca_2501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_806_call_ack_1, ack => zeropad3D_CP_2450_elements(4)); -- 
    rr_2509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(4), ack => type_cast_811_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Sample/ra
      -- 
    ra_2510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_811_inst_ack_0, ack => zeropad3D_CP_2450_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/type_cast_811_Update/ca
      -- 
    ca_2515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_811_inst_ack_1, ack => zeropad3D_CP_2450_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_update_start_
      -- CP-element group 7: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Update/req
      -- 
    ack_2524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_813_inst_ack_0, ack => zeropad3D_CP_2450_elements(7)); -- 
    req_2528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(7), ack => WPIPE_Block0_starting_813_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block0_starting_813_Update/ack
      -- 
    ack_2529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_813_inst_ack_1, ack => zeropad3D_CP_2450_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_update_start_
      -- CP-element group 9: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Update/req
      -- 
    ack_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_816_inst_ack_0, ack => zeropad3D_CP_2450_elements(9)); -- 
    req_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(9), ack => WPIPE_Block1_starting_816_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block1_starting_816_Update/ack
      -- 
    ack_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_816_inst_ack_1, ack => zeropad3D_CP_2450_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_update_start_
      -- CP-element group 11: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Sample/ack
      -- CP-element group 11: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Update/req
      -- 
    ack_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_819_inst_ack_0, ack => zeropad3D_CP_2450_elements(11)); -- 
    req_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(11), ack => WPIPE_Block2_starting_819_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	23 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block2_starting_819_Update/ack
      -- 
    ack_2557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_819_inst_ack_1, ack => zeropad3D_CP_2450_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_update_start_
      -- CP-element group 13: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Sample/ack
      -- CP-element group 13: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Update/req
      -- 
    ack_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_822_inst_ack_0, ack => zeropad3D_CP_2450_elements(13)); -- 
    req_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(13), ack => WPIPE_Block3_starting_822_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	23 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/WPIPE_Block3_starting_822_Update/ack
      -- 
    ack_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_822_inst_ack_1, ack => zeropad3D_CP_2450_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_update_start_
      -- CP-element group 15: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Update/cr
      -- 
    ra_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_826_inst_ack_0, ack => zeropad3D_CP_2450_elements(15)); -- 
    cr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(15), ack => RPIPE_Block0_complete_826_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block0_complete_826_Update/ca
      -- 
    ca_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_826_inst_ack_1, ack => zeropad3D_CP_2450_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_update_start_
      -- CP-element group 17: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Update/cr
      -- 
    ra_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_complete_829_inst_ack_0, ack => zeropad3D_CP_2450_elements(17)); -- 
    cr_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(17), ack => RPIPE_Block1_complete_829_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block1_complete_829_Update/ca
      -- 
    ca_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_complete_829_inst_ack_1, ack => zeropad3D_CP_2450_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_update_start_
      -- CP-element group 19: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Update/cr
      -- 
    ra_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_complete_832_inst_ack_0, ack => zeropad3D_CP_2450_elements(19)); -- 
    cr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(19), ack => RPIPE_Block2_complete_832_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	23 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block2_complete_832_Update/ca
      -- 
    ca_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_complete_832_inst_ack_1, ack => zeropad3D_CP_2450_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_update_start_
      -- CP-element group 21: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Update/cr
      -- 
    ra_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_complete_835_inst_ack_0, ack => zeropad3D_CP_2450_elements(21)); -- 
    cr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(21), ack => RPIPE_Block3_complete_835_inst_req_1); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/RPIPE_Block3_complete_835_Update/ca
      -- 
    ca_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_complete_835_inst_ack_1, ack => zeropad3D_CP_2450_elements(22)); -- 
    -- CP-element group 23:  join  fork  transition  place  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	12 
    -- CP-element group 23: 	14 
    -- CP-element group 23: 	16 
    -- CP-element group 23: 	18 
    -- CP-element group 23: 	20 
    -- CP-element group 23: 	10 
    -- CP-element group 23: 	6 
    -- CP-element group 23: 	8 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	27 
    -- CP-element group 23:  members (13) 
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836__exit__
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_806_to_assign_stmt_836/$exit
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852__entry__
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/$entry
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_update_start_
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Sample/crr
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Update/ccr
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_update_start_
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Update/cr
      -- 
    crr_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(23), ack => call_stmt_839_call_req_0); -- 
    ccr_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(23), ack => call_stmt_839_call_req_1); -- 
    cr_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(23), ack => type_cast_843_inst_req_1); -- 
    zeropad3D_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_2450_elements(12) & zeropad3D_CP_2450_elements(14) & zeropad3D_CP_2450_elements(16) & zeropad3D_CP_2450_elements(18) & zeropad3D_CP_2450_elements(20) & zeropad3D_CP_2450_elements(10) & zeropad3D_CP_2450_elements(6) & zeropad3D_CP_2450_elements(8) & zeropad3D_CP_2450_elements(22);
      gj_zeropad3D_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2450_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Sample/cra
      -- 
    cra_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_839_call_ack_0, ack => zeropad3D_CP_2450_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/call_stmt_839_Update/cca
      -- CP-element group 25: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Sample/rr
      -- 
    cca_2644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_839_call_ack_1, ack => zeropad3D_CP_2450_elements(25)); -- 
    rr_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(25), ack => type_cast_843_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Sample/ra
      -- 
    ra_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_0, ack => zeropad3D_CP_2450_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/type_cast_843_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Sample/req
      -- 
    ca_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_1, ack => zeropad3D_CP_2450_elements(27)); -- 
    req_2666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(27), ack => WPIPE_elapsed_time_pipe_850_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_update_start_
      -- CP-element group 28: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Update/req
      -- 
    ack_2667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_850_inst_ack_0, ack => zeropad3D_CP_2450_elements(28)); -- 
    req_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(28), ack => WPIPE_elapsed_time_pipe_850_inst_req_1); -- 
    -- CP-element group 29:  fork  transition  place  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (13) 
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852__exit__
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854__entry__
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/$exit
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_839_to_assign_stmt_852/WPIPE_elapsed_time_pipe_850_Update/ack
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/$entry
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_update_start_
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Sample/crr
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Update/ccr
      -- 
    ack_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_850_inst_ack_1, ack => zeropad3D_CP_2450_elements(29)); -- 
    crr_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(29), ack => call_stmt_854_call_req_0); -- 
    ccr_2688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2450_elements(29), ack => call_stmt_854_call_req_1); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Sample/cra
      -- 
    cra_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_854_call_ack_0, ack => zeropad3D_CP_2450_elements(30)); -- 
    -- CP-element group 31:  transition  place  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (16) 
      -- CP-element group 31: 	 $exit
      -- CP-element group 31: 	 branch_block_stmt_801/call_stmt_854__exit__
      -- CP-element group 31: 	 branch_block_stmt_801/$exit
      -- CP-element group 31: 	 branch_block_stmt_801/branch_block_stmt_801__exit__
      -- CP-element group 31: 	 branch_block_stmt_801/return__
      -- CP-element group 31: 	 branch_block_stmt_801/merge_stmt_856__exit__
      -- CP-element group 31: 	 branch_block_stmt_801/call_stmt_854/$exit
      -- CP-element group 31: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_801/call_stmt_854/call_stmt_854_Update/cca
      -- CP-element group 31: 	 branch_block_stmt_801/return___PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_801/return___PhiReq/$exit
      -- CP-element group 31: 	 branch_block_stmt_801/merge_stmt_856_PhiReqMerge
      -- CP-element group 31: 	 branch_block_stmt_801/merge_stmt_856_PhiAck/$entry
      -- CP-element group 31: 	 branch_block_stmt_801/merge_stmt_856_PhiAck/$exit
      -- CP-element group 31: 	 branch_block_stmt_801/merge_stmt_856_PhiAck/dummy
      -- 
    cca_2689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_854_call_ack_1, ack => zeropad3D_CP_2450_elements(31)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call10_833 : std_logic_vector(15 downto 0);
    signal call12_836 : std_logic_vector(15 downto 0);
    signal call14_839 : std_logic_vector(63 downto 0);
    signal call1_806 : std_logic_vector(63 downto 0);
    signal call6_827 : std_logic_vector(15 downto 0);
    signal call8_830 : std_logic_vector(15 downto 0);
    signal call_803 : std_logic_vector(15 downto 0);
    signal conv15_844 : std_logic_vector(63 downto 0);
    signal conv_812 : std_logic_vector(63 downto 0);
    signal sub_849 : std_logic_vector(63 downto 0);
    signal type_cast_810_wire : std_logic_vector(63 downto 0);
    signal type_cast_842_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    type_cast_811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_811_inst_req_0;
      type_cast_811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_811_inst_req_1;
      type_cast_811_inst_ack_1<= rack(0);
      type_cast_811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_810_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_812,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_843_inst_req_0;
      type_cast_843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_843_inst_req_1;
      type_cast_843_inst_ack_1<= rack(0);
      type_cast_843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_842_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator SUB_u64_u64_848_inst
    process(conv15_844, conv_812) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv15_844, conv_812, tmp_var);
      sub_849 <= tmp_var; --
    end process;
    -- unary operator type_cast_810_inst
    process(call1_806) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call1_806, tmp_var);
      type_cast_810_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_842_inst
    process(call14_839) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call14_839, tmp_var);
      type_cast_842_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_Block0_complete_826_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_complete_826_inst_req_0;
      RPIPE_Block0_complete_826_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_complete_826_inst_req_1;
      RPIPE_Block0_complete_826_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call6_827 <= data_out(15 downto 0);
      Block0_complete_read_0_gI: SplitGuardInterface generic map(name => "Block0_complete_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_complete_read_0: InputPortRevised -- 
        generic map ( name => "Block0_complete_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_complete_pipe_read_req(0),
          oack => Block0_complete_pipe_read_ack(0),
          odata => Block0_complete_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_complete_829_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_complete_829_inst_req_0;
      RPIPE_Block1_complete_829_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_complete_829_inst_req_1;
      RPIPE_Block1_complete_829_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call8_830 <= data_out(15 downto 0);
      Block1_complete_read_1_gI: SplitGuardInterface generic map(name => "Block1_complete_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_complete_read_1: InputPortRevised -- 
        generic map ( name => "Block1_complete_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_complete_pipe_read_req(0),
          oack => Block1_complete_pipe_read_ack(0),
          odata => Block1_complete_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_complete_832_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_complete_832_inst_req_0;
      RPIPE_Block2_complete_832_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_complete_832_inst_req_1;
      RPIPE_Block2_complete_832_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call10_833 <= data_out(15 downto 0);
      Block2_complete_read_2_gI: SplitGuardInterface generic map(name => "Block2_complete_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_complete_read_2: InputPortRevised -- 
        generic map ( name => "Block2_complete_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_complete_pipe_read_req(0),
          oack => Block2_complete_pipe_read_ack(0),
          odata => Block2_complete_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_complete_835_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_complete_835_inst_req_0;
      RPIPE_Block3_complete_835_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_complete_835_inst_req_1;
      RPIPE_Block3_complete_835_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call12_836 <= data_out(15 downto 0);
      Block3_complete_read_3_gI: SplitGuardInterface generic map(name => "Block3_complete_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_complete_read_3: InputPortRevised -- 
        generic map ( name => "Block3_complete_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_complete_pipe_read_req(0),
          oack => Block3_complete_pipe_read_ack(0),
          odata => Block3_complete_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_starting_813_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_starting_813_inst_req_0;
      WPIPE_Block0_starting_813_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_starting_813_inst_req_1;
      WPIPE_Block0_starting_813_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_803;
      Block0_starting_write_0_gI: SplitGuardInterface generic map(name => "Block0_starting_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_starting_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_starting", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_starting_pipe_write_req(0),
          oack => Block0_starting_pipe_write_ack(0),
          odata => Block0_starting_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_starting_816_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_starting_816_inst_req_0;
      WPIPE_Block1_starting_816_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_starting_816_inst_req_1;
      WPIPE_Block1_starting_816_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_803;
      Block1_starting_write_1_gI: SplitGuardInterface generic map(name => "Block1_starting_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_starting_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_starting", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_starting_pipe_write_req(0),
          oack => Block1_starting_pipe_write_ack(0),
          odata => Block1_starting_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_starting_819_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_starting_819_inst_req_0;
      WPIPE_Block2_starting_819_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_starting_819_inst_req_1;
      WPIPE_Block2_starting_819_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_803;
      Block2_starting_write_2_gI: SplitGuardInterface generic map(name => "Block2_starting_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_starting_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_starting", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_starting_pipe_write_req(0),
          oack => Block2_starting_pipe_write_ack(0),
          odata => Block2_starting_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_starting_822_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_starting_822_inst_req_0;
      WPIPE_Block3_starting_822_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_starting_822_inst_req_1;
      WPIPE_Block3_starting_822_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_803;
      Block3_starting_write_3_gI: SplitGuardInterface generic map(name => "Block3_starting_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_starting_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_starting", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_starting_pipe_write_req(0),
          oack => Block3_starting_pipe_write_ack(0),
          odata => Block3_starting_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_elapsed_time_pipe_850_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_850_inst_req_0;
      WPIPE_elapsed_time_pipe_850_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_850_inst_req_1;
      WPIPE_elapsed_time_pipe_850_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_849;
      elapsed_time_pipe_write_4_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_803_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_803_call_req_0;
      call_stmt_803_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_803_call_req_1;
      call_stmt_803_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_803 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_806_call call_stmt_839_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_806_call_req_0;
      reqL_unguarded(0) <= call_stmt_839_call_req_0;
      call_stmt_806_call_ack_0 <= ackL_unguarded(1);
      call_stmt_839_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_806_call_req_1;
      reqR_unguarded(0) <= call_stmt_839_call_req_1;
      call_stmt_806_call_ack_1 <= ackR_unguarded(1);
      call_stmt_839_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call1_806 <= data_out(127 downto 64);
      call14_839 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_854_call 
    sendOutput_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_854_call_req_0;
      call_stmt_854_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_854_call_req_1;
      call_stmt_854_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_2_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_A is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_A;
architecture zeropad3D_A_arch of zeropad3D_A is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_A_CP_2698_start: Boolean;
  signal zeropad3D_A_CP_2698_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_902_load_0_req_1 : boolean;
  signal ptr_deref_902_load_0_ack_1 : boolean;
  signal ptr_deref_914_load_0_ack_1 : boolean;
  signal type_cast_1467_inst_ack_1 : boolean;
  signal type_cast_1455_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_1 : boolean;
  signal type_cast_969_inst_ack_1 : boolean;
  signal type_cast_1054_inst_ack_0 : boolean;
  signal if_stmt_1063_branch_ack_1 : boolean;
  signal if_stmt_1063_branch_ack_0 : boolean;
  signal phi_stmt_1464_req_0 : boolean;
  signal if_stmt_1063_branch_req_0 : boolean;
  signal phi_stmt_1029_req_0 : boolean;
  signal ptr_deref_1080_load_0_req_1 : boolean;
  signal type_cast_1042_inst_ack_1 : boolean;
  signal ptr_deref_1080_load_0_ack_1 : boolean;
  signal type_cast_1467_inst_req_1 : boolean;
  signal type_cast_1042_inst_req_1 : boolean;
  signal type_cast_969_inst_req_0 : boolean;
  signal type_cast_969_inst_ack_0 : boolean;
  signal type_cast_1054_inst_req_0 : boolean;
  signal ptr_deref_1080_load_0_req_0 : boolean;
  signal phi_stmt_1036_req_1 : boolean;
  signal ptr_deref_1080_load_0_ack_0 : boolean;
  signal type_cast_1054_inst_ack_1 : boolean;
  signal type_cast_969_inst_req_1 : boolean;
  signal ptr_deref_890_load_0_ack_0 : boolean;
  signal ptr_deref_890_load_0_req_0 : boolean;
  signal ptr_deref_914_load_0_req_1 : boolean;
  signal ptr_deref_902_load_0_ack_0 : boolean;
  signal ptr_deref_902_load_0_req_0 : boolean;
  signal ptr_deref_890_load_0_ack_1 : boolean;
  signal ptr_deref_914_load_0_ack_0 : boolean;
  signal ptr_deref_890_load_0_req_1 : boolean;
  signal ptr_deref_914_load_0_req_0 : boolean;
  signal if_stmt_1445_branch_req_0 : boolean;
  signal type_cast_1049_inst_req_0 : boolean;
  signal phi_stmt_1452_ack_0 : boolean;
  signal phi_stmt_1458_ack_0 : boolean;
  signal type_cast_1049_inst_ack_0 : boolean;
  signal type_cast_1049_inst_req_1 : boolean;
  signal type_cast_1049_inst_ack_1 : boolean;
  signal phi_stmt_1043_req_1 : boolean;
  signal if_stmt_1445_branch_ack_1 : boolean;
  signal if_stmt_1445_branch_ack_0 : boolean;
  signal phi_stmt_1029_ack_0 : boolean;
  signal phi_stmt_1036_ack_0 : boolean;
  signal phi_stmt_1043_ack_0 : boolean;
  signal phi_stmt_1464_ack_0 : boolean;
  signal type_cast_1455_inst_ack_1 : boolean;
  signal phi_stmt_1452_req_0 : boolean;
  signal RPIPE_Block0_starting_862_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_862_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_862_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_862_inst_ack_1 : boolean;
  signal LOAD_pad_866_load_0_req_0 : boolean;
  signal LOAD_pad_866_load_0_ack_0 : boolean;
  signal LOAD_pad_866_load_0_req_1 : boolean;
  signal LOAD_pad_866_load_0_ack_1 : boolean;
  signal ptr_deref_878_load_0_req_0 : boolean;
  signal ptr_deref_878_load_0_ack_0 : boolean;
  signal ptr_deref_878_load_0_req_1 : boolean;
  signal ptr_deref_878_load_0_ack_1 : boolean;
  signal if_stmt_1098_branch_req_0 : boolean;
  signal if_stmt_1098_branch_ack_1 : boolean;
  signal if_stmt_1098_branch_ack_0 : boolean;
  signal type_cast_1108_inst_req_0 : boolean;
  signal type_cast_1108_inst_ack_0 : boolean;
  signal type_cast_1108_inst_req_1 : boolean;
  signal type_cast_1108_inst_ack_1 : boolean;
  signal if_stmt_1117_branch_req_0 : boolean;
  signal if_stmt_1117_branch_ack_1 : boolean;
  signal if_stmt_1117_branch_ack_0 : boolean;
  signal ptr_deref_1134_load_0_req_0 : boolean;
  signal ptr_deref_1134_load_0_ack_0 : boolean;
  signal ptr_deref_1134_load_0_req_1 : boolean;
  signal ptr_deref_1134_load_0_ack_1 : boolean;
  signal if_stmt_1152_branch_req_0 : boolean;
  signal if_stmt_1152_branch_ack_1 : boolean;
  signal if_stmt_1152_branch_ack_0 : boolean;
  signal type_cast_1162_inst_req_0 : boolean;
  signal type_cast_1162_inst_ack_0 : boolean;
  signal type_cast_1162_inst_req_1 : boolean;
  signal type_cast_1162_inst_ack_1 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal type_cast_1201_inst_req_0 : boolean;
  signal type_cast_1201_inst_ack_0 : boolean;
  signal type_cast_1201_inst_req_1 : boolean;
  signal type_cast_1201_inst_ack_1 : boolean;
  signal array_obj_ref_1207_index_offset_req_0 : boolean;
  signal array_obj_ref_1207_index_offset_ack_0 : boolean;
  signal array_obj_ref_1207_index_offset_req_1 : boolean;
  signal array_obj_ref_1207_index_offset_ack_1 : boolean;
  signal addr_of_1208_final_reg_req_0 : boolean;
  signal addr_of_1208_final_reg_ack_0 : boolean;
  signal addr_of_1208_final_reg_req_1 : boolean;
  signal addr_of_1208_final_reg_ack_1 : boolean;
  signal ptr_deref_1211_store_0_req_0 : boolean;
  signal ptr_deref_1211_store_0_ack_0 : boolean;
  signal ptr_deref_1211_store_0_req_1 : boolean;
  signal ptr_deref_1211_store_0_ack_1 : boolean;
  signal type_cast_1042_inst_ack_0 : boolean;
  signal type_cast_1042_inst_req_0 : boolean;
  signal type_cast_1220_inst_req_0 : boolean;
  signal type_cast_1220_inst_ack_0 : boolean;
  signal type_cast_1220_inst_req_1 : boolean;
  signal type_cast_1220_inst_ack_1 : boolean;
  signal ptr_deref_1427_load_0_ack_0 : boolean;
  signal ptr_deref_1427_load_0_req_0 : boolean;
  signal type_cast_1467_inst_ack_0 : boolean;
  signal type_cast_1284_inst_req_0 : boolean;
  signal type_cast_1284_inst_ack_0 : boolean;
  signal type_cast_1467_inst_req_0 : boolean;
  signal type_cast_1284_inst_req_1 : boolean;
  signal type_cast_1284_inst_ack_1 : boolean;
  signal phi_stmt_1464_req_1 : boolean;
  signal array_obj_ref_1290_index_offset_req_0 : boolean;
  signal array_obj_ref_1290_index_offset_ack_0 : boolean;
  signal array_obj_ref_1290_index_offset_req_1 : boolean;
  signal array_obj_ref_1290_index_offset_ack_1 : boolean;
  signal addr_of_1291_final_reg_req_0 : boolean;
  signal addr_of_1291_final_reg_ack_0 : boolean;
  signal addr_of_1291_final_reg_req_1 : boolean;
  signal addr_of_1291_final_reg_ack_1 : boolean;
  signal phi_stmt_1458_req_1 : boolean;
  signal type_cast_1463_inst_ack_1 : boolean;
  signal ptr_deref_1295_load_0_req_0 : boolean;
  signal phi_stmt_1029_req_1 : boolean;
  signal ptr_deref_1295_load_0_ack_0 : boolean;
  signal ptr_deref_1295_load_0_req_1 : boolean;
  signal type_cast_1035_inst_ack_1 : boolean;
  signal ptr_deref_1295_load_0_ack_1 : boolean;
  signal type_cast_1035_inst_req_1 : boolean;
  signal type_cast_1309_inst_req_0 : boolean;
  signal type_cast_1309_inst_ack_0 : boolean;
  signal type_cast_1309_inst_req_1 : boolean;
  signal type_cast_1309_inst_ack_1 : boolean;
  signal type_cast_1463_inst_req_1 : boolean;
  signal type_cast_1463_inst_ack_0 : boolean;
  signal type_cast_1035_inst_ack_0 : boolean;
  signal type_cast_1463_inst_req_0 : boolean;
  signal type_cast_1035_inst_req_0 : boolean;
  signal array_obj_ref_1315_index_offset_req_0 : boolean;
  signal array_obj_ref_1315_index_offset_ack_0 : boolean;
  signal array_obj_ref_1315_index_offset_req_1 : boolean;
  signal array_obj_ref_1315_index_offset_ack_1 : boolean;
  signal addr_of_1316_final_reg_req_0 : boolean;
  signal addr_of_1316_final_reg_ack_0 : boolean;
  signal addr_of_1316_final_reg_req_1 : boolean;
  signal addr_of_1316_final_reg_ack_1 : boolean;
  signal WPIPE_Block0_complete_1475_inst_ack_1 : boolean;
  signal WPIPE_Block0_complete_1475_inst_req_1 : boolean;
  signal ptr_deref_1319_store_0_req_0 : boolean;
  signal ptr_deref_1319_store_0_ack_0 : boolean;
  signal ptr_deref_1319_store_0_req_1 : boolean;
  signal ptr_deref_1319_store_0_ack_1 : boolean;
  signal phi_stmt_1452_req_1 : boolean;
  signal type_cast_1327_inst_req_0 : boolean;
  signal type_cast_1327_inst_ack_0 : boolean;
  signal phi_stmt_1458_req_0 : boolean;
  signal type_cast_1327_inst_req_1 : boolean;
  signal type_cast_1327_inst_ack_1 : boolean;
  signal type_cast_1455_inst_ack_0 : boolean;
  signal type_cast_1461_inst_ack_1 : boolean;
  signal type_cast_1461_inst_req_1 : boolean;
  signal if_stmt_1342_branch_req_0 : boolean;
  signal if_stmt_1342_branch_ack_1 : boolean;
  signal if_stmt_1342_branch_ack_0 : boolean;
  signal type_cast_1455_inst_req_0 : boolean;
  signal type_cast_1457_inst_ack_1 : boolean;
  signal type_cast_1457_inst_req_1 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1461_inst_ack_0 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal type_cast_1457_inst_ack_0 : boolean;
  signal type_cast_1457_inst_req_0 : boolean;
  signal phi_stmt_1043_req_0 : boolean;
  signal WPIPE_Block0_complete_1475_inst_ack_0 : boolean;
  signal WPIPE_Block0_complete_1475_inst_req_0 : boolean;
  signal ptr_deref_1378_load_0_req_0 : boolean;
  signal ptr_deref_1378_load_0_ack_0 : boolean;
  signal type_cast_1415_inst_ack_1 : boolean;
  signal ptr_deref_1378_load_0_req_1 : boolean;
  signal ptr_deref_1378_load_0_ack_1 : boolean;
  signal type_cast_1461_inst_req_0 : boolean;
  signal ptr_deref_1427_load_0_ack_1 : boolean;
  signal ptr_deref_1427_load_0_req_1 : boolean;
  signal type_cast_1415_inst_req_1 : boolean;
  signal phi_stmt_1036_req_0 : boolean;
  signal type_cast_1398_inst_req_0 : boolean;
  signal type_cast_1398_inst_ack_0 : boolean;
  signal type_cast_1398_inst_req_1 : boolean;
  signal type_cast_1398_inst_ack_1 : boolean;
  signal type_cast_1415_inst_req_0 : boolean;
  signal type_cast_1415_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_A_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_A_CP_2698_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_A_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2698_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2698_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2698_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_A_CP_2698: Block -- control-path 
    signal zeropad3D_A_CP_2698_elements: BooleanArray(132 downto 0);
    -- 
  begin -- 
    zeropad3D_A_CP_2698_elements(0) <= zeropad3D_A_CP_2698_start;
    zeropad3D_A_CP_2698_symbol <= zeropad3D_A_CP_2698_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_860/$entry
      -- CP-element group 0: 	 branch_block_stmt_860/branch_block_stmt_860__entry__
      -- CP-element group 0: 	 branch_block_stmt_860/assign_stmt_863__entry__
      -- CP-element group 0: 	 branch_block_stmt_860/assign_stmt_863/$entry
      -- CP-element group 0: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Sample/rr
      -- 
    rr_2776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(0), ack => RPIPE_Block0_starting_862_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	132 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	97 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	100 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_860/merge_stmt_1451__exit__
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/$entry
      -- CP-element group 1: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/$entry
      -- 
    cr_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(1), ack => type_cast_1042_inst_req_1); -- 
    rr_3938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(1), ack => type_cast_1049_inst_req_0); -- 
    cr_3943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(1), ack => type_cast_1049_inst_req_1); -- 
    rr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(1), ack => type_cast_1042_inst_req_0); -- 
    cr_3897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(1), ack => type_cast_1035_inst_req_1); -- 
    rr_3892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(1), ack => type_cast_1035_inst_req_0); -- 
    zeropad3D_A_CP_2698_elements(1) <= zeropad3D_A_CP_2698_elements(132);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_update_start_
      -- CP-element group 2: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Update/cr
      -- 
    ra_2777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_862_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(2)); -- 
    cr_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(2), ack => RPIPE_Block0_starting_862_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3: 	7 
    -- CP-element group 3: 	11 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	15 
    -- CP-element group 3: 	10 
    -- CP-element group 3: 	9 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (126) 
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_update_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_update_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_update_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_863__exit__
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026__entry__
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_863/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_863/RPIPE_Block0_starting_862_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_update_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_update_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_update_start_
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_base_plus_offset/sum_rename_ack
      -- 
    ca_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_862_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(3)); -- 
    cr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_902_load_0_req_1); -- 
    cr_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => type_cast_969_inst_req_1); -- 
    rr_2901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_890_load_0_req_0); -- 
    cr_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_914_load_0_req_1); -- 
    rr_2951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_902_load_0_req_0); -- 
    cr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_890_load_0_req_1); -- 
    rr_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_914_load_0_req_0); -- 
    rr_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => LOAD_pad_866_load_0_req_0); -- 
    cr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => LOAD_pad_866_load_0_req_1); -- 
    rr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_878_load_0_req_0); -- 
    cr_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(3), ack => ptr_deref_878_load_0_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/word_access_start/$exit
      -- CP-element group 4: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Sample/word_access_start/word_0/ra
      -- 
    ra_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_866_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	14 
    -- CP-element group 5:  members (12) 
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/word_access_complete/word_0/ca
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/LOAD_pad_866_Merge/$entry
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/LOAD_pad_866_Merge/$exit
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/LOAD_pad_866_Merge/merge_req
      -- CP-element group 5: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/LOAD_pad_866_Update/LOAD_pad_866_Merge/merge_ack
      -- 
    ca_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_866_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(5)); -- 
    rr_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(5), ack => type_cast_969_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Sample/word_access_start/word_0/ra
      -- 
    ra_2852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_878_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	3 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/word_access_complete/word_0/ca
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/ptr_deref_878_Merge/$entry
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/ptr_deref_878_Merge/$exit
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/ptr_deref_878_Merge/merge_req
      -- CP-element group 7: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_878_Update/ptr_deref_878_Merge/merge_ack
      -- 
    ca_2863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_878_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_sample_completed_
      -- 
    ra_2902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_890_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	3 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/ptr_deref_890_Merge/merge_ack
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/ptr_deref_890_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/ptr_deref_890_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/ptr_deref_890_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_890_update_completed_
      -- 
    ca_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_890_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/word_access_start/word_0/ra
      -- CP-element group 10: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Sample/word_access_start/$exit
      -- 
    ra_2952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	16 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/word_access_complete/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/word_access_complete/word_0/ca
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/word_access_complete/$exit
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/ptr_deref_902_Merge/$entry
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/ptr_deref_902_Merge/merge_req
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/ptr_deref_902_Merge/$exit
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/ptr_deref_902_Merge/merge_ack
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_902_Update/$exit
      -- 
    ca_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/word_access_start/word_0/ra
      -- CP-element group 12: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Sample/word_access_start/$exit
      -- 
    ra_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_914_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/ptr_deref_914_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/ptr_deref_914_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/ptr_deref_914_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/ptr_deref_914_Merge/merge_ack
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/ptr_deref_914_Update/$exit
      -- 
    ca_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_914_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	5 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Sample/ra
      -- 
    ra_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_969_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/type_cast_969_Update/$exit
      -- 
    ca_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_969_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(15)); -- 
    -- CP-element group 16:  join  fork  transition  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	15 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	89 
    -- CP-element group 16: 	90 
    -- CP-element group 16: 	91 
    -- CP-element group 16:  members (10) 
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1036/$entry
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$entry
      -- CP-element group 16: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026__exit__
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody
      -- CP-element group 16: 	 branch_block_stmt_860/assign_stmt_867_to_assign_stmt_1026/$exit
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/$entry
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1029/$entry
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$entry
      -- CP-element group 16: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1043/$entry
      -- 
    zeropad3D_A_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(7) & zeropad3D_A_CP_2698_elements(11) & zeropad3D_A_CP_2698_elements(15) & zeropad3D_A_CP_2698_elements(9) & zeropad3D_A_CP_2698_elements(13);
      gj_zeropad3D_A_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	107 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Sample/$exit
      -- 
    ra_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(17)); -- 
    -- CP-element group 18:  branch  transition  place  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	107 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (13) 
      -- CP-element group 18: 	 branch_block_stmt_860/R_cmp_1064_place
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063_if_link/$entry
      -- CP-element group 18: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063_else_link/$entry
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063_eval_test/$exit
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063_eval_test/branch_req
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063_dead_link/$entry
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063_eval_test/$entry
      -- CP-element group 18: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/$exit
      -- CP-element group 18: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062__exit__
      -- CP-element group 18: 	 branch_block_stmt_860/if_stmt_1063__entry__
      -- 
    ca_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(18)); -- 
    branch_req_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(18), ack => if_stmt_1063_branch_req_0); -- 
    -- CP-element group 19:  transition  place  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	108 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_860/whilex_xbody_ifx_xthen
      -- CP-element group 19: 	 branch_block_stmt_860/if_stmt_1063_if_link/$exit
      -- CP-element group 19: 	 branch_block_stmt_860/if_stmt_1063_if_link/if_choice_transition
      -- CP-element group 19: 	 branch_block_stmt_860/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 19: 	 branch_block_stmt_860/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- 
    if_choice_transition_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1063_branch_ack_1, ack => zeropad3D_A_CP_2698_elements(19)); -- 
    -- CP-element group 20:  merge  transition  place  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (11) 
      -- CP-element group 20: 	 branch_block_stmt_860/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 20: 	 branch_block_stmt_860/merge_stmt_1069_PhiReqMerge
      -- CP-element group 20: 	 branch_block_stmt_860/if_stmt_1063_else_link/else_choice_transition
      -- CP-element group 20: 	 branch_block_stmt_860/if_stmt_1063_else_link/$exit
      -- CP-element group 20: 	 branch_block_stmt_860/merge_stmt_1069__exit__
      -- CP-element group 20: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097__entry__
      -- CP-element group 20: 	 branch_block_stmt_860/merge_stmt_1069_PhiAck/dummy
      -- CP-element group 20: 	 branch_block_stmt_860/merge_stmt_1069_PhiAck/$exit
      -- CP-element group 20: 	 branch_block_stmt_860/merge_stmt_1069_PhiAck/$entry
      -- CP-element group 20: 	 branch_block_stmt_860/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 20: 	 branch_block_stmt_860/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- 
    else_choice_transition_3066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1063_branch_ack_0, ack => zeropad3D_A_CP_2698_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (27) 
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_update_start_
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/word_access_complete/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/word_access_complete/word_0/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/word_access_complete/word_0/cr
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_addr_resize/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_addr_resize/$exit
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_word_addrgen/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_word_addrgen/$exit
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_word_addrgen/root_register_req
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_word_addrgen/root_register_ack
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_word_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/word_access_start/word_0/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/word_access_start/word_0/rr
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_plus_offset/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_plus_offset/$exit
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/word_access_start/$entry
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_root_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_address_resized
      -- CP-element group 21: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_base_addr_resize/base_resize_req
      -- 
    cr_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(21), ack => ptr_deref_1080_load_0_req_1); -- 
    rr_3104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(21), ack => ptr_deref_1080_load_0_req_0); -- 
    zeropad3D_A_CP_2698_elements(21) <= zeropad3D_A_CP_2698_elements(20);
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/word_access_start/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/word_access_start/word_0/ra
      -- CP-element group 22: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Sample/word_access_start/$exit
      -- 
    ra_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1080_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(22)); -- 
    -- CP-element group 23:  branch  transition  place  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (19) 
      -- CP-element group 23: 	 branch_block_stmt_860/R_cmp45_1099_place
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/word_access_complete/$exit
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/word_access_complete/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/word_access_complete/word_0/ca
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/ptr_deref_1080_Merge/$entry
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/ptr_deref_1080_Merge/$exit
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/ptr_deref_1080_Merge/merge_req
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/ptr_deref_1080_Update/ptr_deref_1080_Merge/merge_ack
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097/$exit
      -- CP-element group 23: 	 branch_block_stmt_860/assign_stmt_1077_to_assign_stmt_1097__exit__
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098__entry__
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098_dead_link/$entry
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098_eval_test/$entry
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098_eval_test/$exit
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098_eval_test/branch_req
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098_if_link/$entry
      -- CP-element group 23: 	 branch_block_stmt_860/if_stmt_1098_else_link/$entry
      -- 
    ca_3116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1080_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(23)); -- 
    branch_req_3129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(23), ack => if_stmt_1098_branch_req_0); -- 
    -- CP-element group 24:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (18) 
      -- CP-element group 24: 	 branch_block_stmt_860/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse47
      -- CP-element group 24: 	 branch_block_stmt_860/merge_stmt_1104_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_860/merge_stmt_1104__exit__
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116__entry__
      -- CP-element group 24: 	 branch_block_stmt_860/if_stmt_1098_if_link/$exit
      -- CP-element group 24: 	 branch_block_stmt_860/if_stmt_1098_if_link/if_choice_transition
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/$entry
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_update_start_
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_860/merge_stmt_1104_PhiAck/dummy
      -- CP-element group 24: 	 branch_block_stmt_860/merge_stmt_1104_PhiAck/$exit
      -- CP-element group 24: 	 branch_block_stmt_860/merge_stmt_1104_PhiAck/$entry
      -- CP-element group 24: 	 branch_block_stmt_860/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse47_PhiReq/$exit
      -- CP-element group 24: 	 branch_block_stmt_860/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse47_PhiReq/$entry
      -- 
    if_choice_transition_3134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1098_branch_ack_1, ack => zeropad3D_A_CP_2698_elements(24)); -- 
    rr_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(24), ack => type_cast_1108_inst_req_0); -- 
    cr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(24), ack => type_cast_1108_inst_req_1); -- 
    -- CP-element group 25:  transition  place  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	108 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_860/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 25: 	 branch_block_stmt_860/if_stmt_1098_else_link/$exit
      -- CP-element group 25: 	 branch_block_stmt_860/if_stmt_1098_else_link/else_choice_transition
      -- CP-element group 25: 	 branch_block_stmt_860/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- CP-element group 25: 	 branch_block_stmt_860/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- 
    else_choice_transition_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1098_branch_ack_0, ack => zeropad3D_A_CP_2698_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Sample/ra
      -- 
    ra_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1108_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(26)); -- 
    -- CP-element group 27:  branch  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (13) 
      -- CP-element group 27: 	 branch_block_stmt_860/R_cmp52_1118_place
      -- CP-element group 27: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116__exit__
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117__entry__
      -- CP-element group 27: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/$exit
      -- CP-element group 27: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_860/assign_stmt_1109_to_assign_stmt_1116/type_cast_1108_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117_dead_link/$entry
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117_eval_test/$entry
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117_eval_test/$exit
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117_eval_test/branch_req
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117_if_link/$entry
      -- CP-element group 27: 	 branch_block_stmt_860/if_stmt_1117_else_link/$entry
      -- 
    ca_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1108_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(27)); -- 
    branch_req_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(27), ack => if_stmt_1117_branch_req_0); -- 
    -- CP-element group 28:  transition  place  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	108 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 branch_block_stmt_860/lorx_xlhsx_xfalse47_ifx_xthen
      -- CP-element group 28: 	 branch_block_stmt_860/lorx_xlhsx_xfalse47_ifx_xthen_PhiReq/$entry
      -- CP-element group 28: 	 branch_block_stmt_860/lorx_xlhsx_xfalse47_ifx_xthen_PhiReq/$exit
      -- CP-element group 28: 	 branch_block_stmt_860/if_stmt_1117_if_link/$exit
      -- CP-element group 28: 	 branch_block_stmt_860/if_stmt_1117_if_link/if_choice_transition
      -- 
    if_choice_transition_3170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1117_branch_ack_1, ack => zeropad3D_A_CP_2698_elements(28)); -- 
    -- CP-element group 29:  merge  transition  place  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (11) 
      -- CP-element group 29: 	 branch_block_stmt_860/lorx_xlhsx_xfalse47_lorx_xlhsx_xfalse54
      -- CP-element group 29: 	 branch_block_stmt_860/merge_stmt_1123_PhiAck/$exit
      -- CP-element group 29: 	 branch_block_stmt_860/merge_stmt_1123_PhiAck/$entry
      -- CP-element group 29: 	 branch_block_stmt_860/merge_stmt_1123_PhiAck/dummy
      -- CP-element group 29: 	 branch_block_stmt_860/merge_stmt_1123_PhiReqMerge
      -- CP-element group 29: 	 branch_block_stmt_860/merge_stmt_1123__exit__
      -- CP-element group 29: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151__entry__
      -- CP-element group 29: 	 branch_block_stmt_860/if_stmt_1117_else_link/$exit
      -- CP-element group 29: 	 branch_block_stmt_860/if_stmt_1117_else_link/else_choice_transition
      -- CP-element group 29: 	 branch_block_stmt_860/lorx_xlhsx_xfalse47_lorx_xlhsx_xfalse54_PhiReq/$exit
      -- CP-element group 29: 	 branch_block_stmt_860/lorx_xlhsx_xfalse47_lorx_xlhsx_xfalse54_PhiReq/$entry
      -- 
    else_choice_transition_3174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1117_branch_ack_0, ack => zeropad3D_A_CP_2698_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (27) 
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_update_start_
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_address_calculated
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_word_address_calculated
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_root_address_calculated
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_address_resized
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_addr_resize/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_addr_resize/$exit
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_addr_resize/base_resize_req
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_addr_resize/base_resize_ack
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_plus_offset/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_plus_offset/$exit
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_word_addrgen/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_word_addrgen/$exit
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_word_addrgen/root_register_req
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_word_addrgen/root_register_ack
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/word_access_start/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/word_access_start/word_0/rr
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/word_access_complete/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/word_access_complete/word_0/$entry
      -- CP-element group 30: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/word_access_complete/word_0/cr
      -- 
    cr_3223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(30), ack => ptr_deref_1134_load_0_req_1); -- 
    rr_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(30), ack => ptr_deref_1134_load_0_req_0); -- 
    zeropad3D_A_CP_2698_elements(30) <= zeropad3D_A_CP_2698_elements(29);
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Sample/word_access_start/word_0/ra
      -- 
    ra_3213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(31)); -- 
    -- CP-element group 32:  branch  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (19) 
      -- CP-element group 32: 	 branch_block_stmt_860/R_cmp62_1153_place
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151__exit__
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152__entry__
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/$exit
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/ptr_deref_1134_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/ptr_deref_1134_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/ptr_deref_1134_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_860/assign_stmt_1131_to_assign_stmt_1151/ptr_deref_1134_Update/ptr_deref_1134_Merge/merge_ack
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152_dead_link/$entry
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152_eval_test/$entry
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152_eval_test/$exit
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152_eval_test/branch_req
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152_if_link/$entry
      -- CP-element group 32: 	 branch_block_stmt_860/if_stmt_1152_else_link/$entry
      -- 
    ca_3224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(32)); -- 
    branch_req_3237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(32), ack => if_stmt_1152_branch_req_0); -- 
    -- CP-element group 33:  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	49 
    -- CP-element group 33: 	50 
    -- CP-element group 33: 	52 
    -- CP-element group 33: 	54 
    -- CP-element group 33: 	56 
    -- CP-element group 33: 	58 
    -- CP-element group 33: 	60 
    -- CP-element group 33: 	62 
    -- CP-element group 33: 	64 
    -- CP-element group 33: 	67 
    -- CP-element group 33:  members (46) 
      -- CP-element group 33: 	 branch_block_stmt_860/lorx_xlhsx_xfalse54_ifx_xelse
      -- CP-element group 33: 	 branch_block_stmt_860/merge_stmt_1216_PhiReqMerge
      -- CP-element group 33: 	 branch_block_stmt_860/merge_stmt_1216__exit__
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321__entry__
      -- CP-element group 33: 	 branch_block_stmt_860/if_stmt_1152_if_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_860/if_stmt_1152_if_link/if_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_update_start
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Update/req
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_complete/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_complete/req
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/word_access_complete/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/word_access_complete/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/word_access_complete/word_0/cr
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_update_start
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Update/req
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_complete/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_complete/req
      -- CP-element group 33: 	 branch_block_stmt_860/merge_stmt_1216_PhiAck/dummy
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_update_start_
      -- CP-element group 33: 	 branch_block_stmt_860/merge_stmt_1216_PhiAck/$exit
      -- CP-element group 33: 	 branch_block_stmt_860/merge_stmt_1216_PhiAck/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/lorx_xlhsx_xfalse54_ifx_xelse_PhiReq/$exit
      -- CP-element group 33: 	 branch_block_stmt_860/lorx_xlhsx_xfalse54_ifx_xelse_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/word_access_complete/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/word_access_complete/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/word_access_complete/word_0/cr
      -- 
    if_choice_transition_3242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1152_branch_ack_1, ack => zeropad3D_A_CP_2698_elements(33)); -- 
    rr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => type_cast_1220_inst_req_0); -- 
    cr_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => type_cast_1220_inst_req_1); -- 
    cr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => type_cast_1284_inst_req_1); -- 
    req_3450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => array_obj_ref_1290_index_offset_req_1); -- 
    req_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => addr_of_1291_final_reg_req_1); -- 
    cr_3510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => ptr_deref_1295_load_0_req_1); -- 
    cr_3529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => type_cast_1309_inst_req_1); -- 
    req_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => array_obj_ref_1315_index_offset_req_1); -- 
    req_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => addr_of_1316_final_reg_req_1); -- 
    cr_3625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(33), ack => ptr_deref_1319_store_0_req_1); -- 
    -- CP-element group 34:  transition  place  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	108 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_860/lorx_xlhsx_xfalse54_ifx_xthen
      -- CP-element group 34: 	 branch_block_stmt_860/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_860/if_stmt_1152_else_link/$exit
      -- CP-element group 34: 	 branch_block_stmt_860/if_stmt_1152_else_link/else_choice_transition
      -- CP-element group 34: 	 branch_block_stmt_860/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1152_branch_ack_0, ack => zeropad3D_A_CP_2698_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	108 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Sample/ra
      -- 
    ra_3260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	108 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	39 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Update/ca
      -- 
    ca_3265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	108 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Sample/ra
      -- 
    ra_3274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	108 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Update/ca
      -- 
    ca_3279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	36 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Sample/rr
      -- 
    rr_3287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(39), ack => type_cast_1201_inst_req_0); -- 
    zeropad3D_A_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(36) & zeropad3D_A_CP_2698_elements(38);
      gj_zeropad3D_A_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Sample/ra
      -- 
    ra_3288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	108 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (16) 
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_resized_1
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_scaled_1
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_computed_1
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_resize_1/$entry
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_resize_1/$exit
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_resize_1/index_resize_req
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_resize_1/index_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_scale_1/$entry
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_scale_1/$exit
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_scale_1/scale_rename_req
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_index_scale_1/scale_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Sample/req
      -- 
    ca_3293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(41)); -- 
    req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(41), ack => array_obj_ref_1207_index_offset_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	48 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_sample_complete
      -- CP-element group 42: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Sample/ack
      -- 
    ack_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1207_index_offset_ack_0, ack => zeropad3D_A_CP_2698_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	108 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (11) 
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_offset_calculated
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Update/ack
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_request/$entry
      -- CP-element group 43: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_request/req
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1207_index_offset_ack_1, ack => zeropad3D_A_CP_2698_elements(43)); -- 
    req_3333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(43), ack => addr_of_1208_final_reg_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_request/$exit
      -- CP-element group 44: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_request/ack
      -- 
    ack_3334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1208_final_reg_ack_0, ack => zeropad3D_A_CP_2698_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	108 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (28) 
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_complete/ack
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_word_addrgen/root_register_ack
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/ptr_deref_1211_Split/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/ptr_deref_1211_Split/$exit
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/ptr_deref_1211_Split/split_req
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/ptr_deref_1211_Split/split_ack
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/word_access_start/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/word_access_start/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/word_access_start/word_0/rr
      -- 
    ack_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1208_final_reg_ack_1, ack => zeropad3D_A_CP_2698_elements(45)); -- 
    rr_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(45), ack => ptr_deref_1211_store_0_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/word_access_start/$exit
      -- CP-element group 46: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Sample/word_access_start/word_0/ra
      -- 
    ra_3378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1211_store_0_ack_0, ack => zeropad3D_A_CP_2698_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	108 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/word_access_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/word_access_complete/word_0/ca
      -- 
    ca_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1211_store_0_ack_1, ack => zeropad3D_A_CP_2698_elements(47)); -- 
    -- CP-element group 48:  join  transition  place  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	42 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	109 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214__exit__
      -- CP-element group 48: 	 branch_block_stmt_860/ifx_xthen_ifx_xend
      -- CP-element group 48: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/$exit
      -- CP-element group 48: 	 branch_block_stmt_860/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_860/ifx_xthen_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_A_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(42) & zeropad3D_A_CP_2698_elements(47);
      gj_zeropad3D_A_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	33 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Sample/ra
      -- 
    ra_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	33 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	59 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1220_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Sample/rr
      -- 
    ca_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(50)); -- 
    rr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(50), ack => type_cast_1284_inst_req_0); -- 
    rr_3524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(50), ack => type_cast_1309_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Sample/ra
      -- 
    ra_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	33 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (16) 
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1284_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_resized_1
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_scaled_1
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_computed_1
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_resize_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_resize_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_resize_1/index_resize_req
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_resize_1/index_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_scale_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_scale_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_scale_1/scale_rename_req
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_index_scale_1/scale_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Sample/req
      -- 
    ca_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(52)); -- 
    req_3445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(52), ack => array_obj_ref_1290_index_offset_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	68 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_sample_complete
      -- CP-element group 53: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Sample/ack
      -- 
    ack_3446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1290_index_offset_ack_0, ack => zeropad3D_A_CP_2698_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	33 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (11) 
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_root_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_offset_calculated
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_final_index_sum_regn_Update/ack
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_base_plus_offset/$entry
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_base_plus_offset/$exit
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1290_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_request/$entry
      -- CP-element group 54: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_request/req
      -- 
    ack_3451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1290_index_offset_ack_1, ack => zeropad3D_A_CP_2698_elements(54)); -- 
    req_3460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(54), ack => addr_of_1291_final_reg_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_request/$exit
      -- CP-element group 55: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_request/ack
      -- 
    ack_3461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1291_final_reg_ack_0, ack => zeropad3D_A_CP_2698_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	33 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_complete/$exit
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1291_complete/ack
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/word_access_start/word_0/rr
      -- 
    ack_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1291_final_reg_ack_1, ack => zeropad3D_A_CP_2698_elements(56)); -- 
    rr_3499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(56), ack => ptr_deref_1295_load_0_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/word_access_start/$exit
      -- CP-element group 57: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/word_access_start/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Sample/word_access_start/word_0/ra
      -- 
    ra_3500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1295_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	33 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	65 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/word_access_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/word_access_complete/word_0/$exit
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/word_access_complete/word_0/ca
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/ptr_deref_1295_Merge/$entry
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/ptr_deref_1295_Merge/$exit
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/ptr_deref_1295_Merge/merge_req
      -- CP-element group 58: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1295_Update/ptr_deref_1295_Merge/merge_ack
      -- 
    ca_3511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1295_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	50 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Sample/ra
      -- 
    ra_3525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1309_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	33 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (16) 
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/type_cast_1309_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_scale_1/scale_rename_req
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Sample/req
      -- 
    ca_3530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1309_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(60)); -- 
    req_3555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(60), ack => array_obj_ref_1315_index_offset_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	68 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Sample/ack
      -- 
    ack_3556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1315_index_offset_ack_0, ack => zeropad3D_A_CP_2698_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	33 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (11) 
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_offset_calculated
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_final_index_sum_regn_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/array_obj_ref_1315_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_request/$entry
      -- CP-element group 62: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_request/req
      -- 
    ack_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1315_index_offset_ack_1, ack => zeropad3D_A_CP_2698_elements(62)); -- 
    req_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(62), ack => addr_of_1316_final_reg_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_request/$exit
      -- CP-element group 63: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_request/ack
      -- 
    ack_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1316_final_reg_ack_0, ack => zeropad3D_A_CP_2698_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	33 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (19) 
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/addr_of_1316_complete/ack
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_word_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_address_resized
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_addr_resize/$entry
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_addr_resize/$exit
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_addr_resize/base_resize_req
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_addr_resize/base_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_word_addrgen/$entry
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_word_addrgen/$exit
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_word_addrgen/root_register_req
      -- CP-element group 64: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_word_addrgen/root_register_ack
      -- 
    ack_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1316_final_reg_ack_1, ack => zeropad3D_A_CP_2698_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	58 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (9) 
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/ptr_deref_1319_Split/$entry
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/ptr_deref_1319_Split/$exit
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/ptr_deref_1319_Split/split_req
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/ptr_deref_1319_Split/split_ack
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/word_access_start/$entry
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/word_access_start/word_0/$entry
      -- CP-element group 65: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/word_access_start/word_0/rr
      -- 
    rr_3614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(65), ack => ptr_deref_1319_store_0_req_0); -- 
    zeropad3D_A_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(58) & zeropad3D_A_CP_2698_elements(64);
      gj_zeropad3D_A_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/word_access_start/$exit
      -- CP-element group 66: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/word_access_start/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Sample/word_access_start/word_0/ra
      -- 
    ra_3615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1319_store_0_ack_0, ack => zeropad3D_A_CP_2698_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	33 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (5) 
      -- CP-element group 67: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/word_access_complete/$exit
      -- CP-element group 67: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/word_access_complete/word_0/$exit
      -- CP-element group 67: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/ptr_deref_1319_Update/word_access_complete/word_0/ca
      -- 
    ca_3626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1319_store_0_ack_1, ack => zeropad3D_A_CP_2698_elements(67)); -- 
    -- CP-element group 68:  join  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	53 
    -- CP-element group 68: 	61 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	109 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321__exit__
      -- CP-element group 68: 	 branch_block_stmt_860/ifx_xelse_ifx_xend
      -- CP-element group 68: 	 branch_block_stmt_860/assign_stmt_1221_to_assign_stmt_1321/$exit
      -- CP-element group 68: 	 branch_block_stmt_860/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_860/ifx_xelse_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_A_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(53) & zeropad3D_A_CP_2698_elements(61) & zeropad3D_A_CP_2698_elements(67);
      gj_zeropad3D_A_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	109 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Sample/ra
      -- 
    ra_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1327_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	109 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341__exit__
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342__entry__
      -- CP-element group 70: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/$exit
      -- CP-element group 70: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_860/R_cmp131_1343_place
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_860/if_stmt_1342_else_link/$entry
      -- 
    ca_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1327_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(70)); -- 
    branch_req_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(70), ack => if_stmt_1342_branch_req_0); -- 
    -- CP-element group 71:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71: 	119 
    -- CP-element group 71: 	121 
    -- CP-element group 71: 	122 
    -- CP-element group 71: 	124 
    -- CP-element group 71: 	125 
    -- CP-element group 71:  members (40) 
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Update/cr
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/cr
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/merge_stmt_1348_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_860/merge_stmt_1348__exit__
      -- CP-element group 71: 	 branch_block_stmt_860/assign_stmt_1354__entry__
      -- CP-element group 71: 	 branch_block_stmt_860/assign_stmt_1354__exit__
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/merge_stmt_1348_PhiAck/dummy
      -- CP-element group 71: 	 branch_block_stmt_860/merge_stmt_1348_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/merge_stmt_1348_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xend_ifx_xthen133_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xend_ifx_xthen133_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Update/cr
      -- CP-element group 71: 	 branch_block_stmt_860/if_stmt_1342_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_860/if_stmt_1342_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xend_ifx_xthen133
      -- CP-element group 71: 	 branch_block_stmt_860/assign_stmt_1354/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/assign_stmt_1354/$exit
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Sample/rr
      -- 
    if_choice_transition_3656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1342_branch_ack_1, ack => zeropad3D_A_CP_2698_elements(71)); -- 
    cr_4133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(71), ack => type_cast_1455_inst_req_1); -- 
    cr_4179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(71), ack => type_cast_1467_inst_req_1); -- 
    rr_4174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(71), ack => type_cast_1467_inst_req_0); -- 
    cr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(71), ack => type_cast_1461_inst_req_1); -- 
    rr_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(71), ack => type_cast_1455_inst_req_0); -- 
    rr_4151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(71), ack => type_cast_1461_inst_req_0); -- 
    -- CP-element group 72:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	75 
    -- CP-element group 72: 	76 
    -- CP-element group 72: 	79 
    -- CP-element group 72: 	81 
    -- CP-element group 72: 	82 
    -- CP-element group 72: 	83 
    -- CP-element group 72:  members (76) 
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/word_access_complete/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/merge_stmt_1356_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/merge_stmt_1356_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_860/merge_stmt_1356_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/word_access_complete/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_860/merge_stmt_1356__exit__
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444__entry__
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/merge_stmt_1356_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/word_access_start/word_0/rr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_update_start_
      -- CP-element group 72: 	 branch_block_stmt_860/ifx_xend_ifx_xelse138_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/ifx_xend_ifx_xelse138_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/word_access_start/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_word_addrgen/root_register_ack
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_860/if_stmt_1342_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/if_stmt_1342_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/ifx_xend_ifx_xelse138
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_update_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_update_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_word_addrgen/root_register_ack
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/word_access_start/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/word_access_start/word_0/rr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/word_access_complete/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/word_access_complete/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/word_access_complete/word_0/cr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/word_access_complete/word_0/cr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_update_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_update_start_
      -- CP-element group 72: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Update/$entry
      -- 
    else_choice_transition_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1342_branch_ack_0, ack => zeropad3D_A_CP_2698_elements(72)); -- 
    rr_3793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => ptr_deref_1427_load_0_req_0); -- 
    rr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => type_cast_1366_inst_req_0); -- 
    cr_3681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => type_cast_1366_inst_req_1); -- 
    rr_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => ptr_deref_1378_load_0_req_0); -- 
    cr_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => ptr_deref_1378_load_0_req_1); -- 
    cr_3804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => ptr_deref_1427_load_0_req_1); -- 
    cr_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => type_cast_1415_inst_req_1); -- 
    cr_3745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(72), ack => type_cast_1398_inst_req_1); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Sample/ra
      -- 
    ra_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	77 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1366_Update/ca
      -- 
    ca_3682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/word_access_start/$exit
      -- CP-element group 75: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/word_access_start/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Sample/word_access_start/word_0/ra
      -- 
    ra_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1378_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	72 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/word_access_complete/$exit
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/word_access_complete/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/word_access_complete/word_0/ca
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/ptr_deref_1378_Merge/$entry
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/ptr_deref_1378_Merge/$exit
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/ptr_deref_1378_Merge/merge_req
      -- CP-element group 76: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1378_Update/ptr_deref_1378_Merge/merge_ack
      -- 
    ca_3727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1378_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Sample/rr
      -- 
    rr_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(77), ack => type_cast_1398_inst_req_0); -- 
    zeropad3D_A_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(74) & zeropad3D_A_CP_2698_elements(76);
      gj_zeropad3D_A_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Sample/ra
      -- 
    ra_3741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(78)); -- 
    -- CP-element group 79:  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	72 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1398_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Sample/rr
      -- 
    ca_3746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(79)); -- 
    rr_3754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(79), ack => type_cast_1415_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Sample/ra
      -- 
    ra_3755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	72 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	84 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/type_cast_1415_Update/$exit
      -- 
    ca_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/word_access_start/word_0/ra
      -- CP-element group 82: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/word_access_start/$exit
      -- CP-element group 82: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Sample/$exit
      -- 
    ra_3794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1427_load_0_ack_0, ack => zeropad3D_A_CP_2698_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	72 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/word_access_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/ptr_deref_1427_Merge/merge_ack
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/ptr_deref_1427_Merge/$exit
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/ptr_deref_1427_Merge/merge_req
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/ptr_deref_1427_Merge/$entry
      -- CP-element group 83: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/ptr_deref_1427_Update/word_access_complete/word_0/ca
      -- 
    ca_3805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1427_load_0_ack_1, ack => zeropad3D_A_CP_2698_elements(83)); -- 
    -- CP-element group 84:  branch  join  transition  place  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	81 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (10) 
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445_else_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444__exit__
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445__entry__
      -- CP-element group 84: 	 branch_block_stmt_860/if_stmt_1445_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_860/assign_stmt_1362_to_assign_stmt_1444/$exit
      -- CP-element group 84: 	 branch_block_stmt_860/R_cmp162_1446_place
      -- 
    branch_req_3818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(84), ack => if_stmt_1445_branch_req_0); -- 
    zeropad3D_A_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(81) & zeropad3D_A_CP_2698_elements(83);
      gj_zeropad3D_A_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_860/if_stmt_1445_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_860/if_stmt_1445_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_860/ifx_xelse138_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_860/assign_stmt_1477/$entry
      -- CP-element group 85: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_860/ifx_xelse138_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_860/merge_stmt_1473__exit__
      -- CP-element group 85: 	 branch_block_stmt_860/assign_stmt_1477__entry__
      -- CP-element group 85: 	 branch_block_stmt_860/ifx_xelse138_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_860/merge_stmt_1473_PhiAck/dummy
      -- CP-element group 85: 	 branch_block_stmt_860/merge_stmt_1473_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_860/merge_stmt_1473_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_860/merge_stmt_1473_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Sample/req
      -- 
    if_choice_transition_3823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1445_branch_ack_1, ack => zeropad3D_A_CP_2698_elements(85)); -- 
    req_3840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(85), ack => WPIPE_Block0_complete_1475_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	110 
    -- CP-element group 86: 	111 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	114 
    -- CP-element group 86: 	116 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/if_stmt_1445_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_860/if_stmt_1445_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1464/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/$entry
      -- 
    else_choice_transition_3827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1445_branch_ack_0, ack => zeropad3D_A_CP_2698_elements(86)); -- 
    cr_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(86), ack => type_cast_1463_inst_req_1); -- 
    rr_4094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(86), ack => type_cast_1463_inst_req_0); -- 
    cr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(86), ack => type_cast_1457_inst_req_1); -- 
    rr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(86), ack => type_cast_1457_inst_req_0); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_update_start_
      -- CP-element group 87: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Update/req
      -- CP-element group 87: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Sample/$exit
      -- 
    ack_3841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1475_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(87)); -- 
    req_3845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(87), ack => WPIPE_Block0_complete_1475_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_860/assign_stmt_1477/$exit
      -- CP-element group 88: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_update_completed_
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_860/$exit
      -- CP-element group 88: 	 branch_block_stmt_860/branch_block_stmt_860__exit__
      -- CP-element group 88: 	 branch_block_stmt_860/assign_stmt_1477__exit__
      -- CP-element group 88: 	 branch_block_stmt_860/return__
      -- CP-element group 88: 	 branch_block_stmt_860/merge_stmt_1479__exit__
      -- CP-element group 88: 	 branch_block_stmt_860/merge_stmt_1479_PhiAck/dummy
      -- CP-element group 88: 	 branch_block_stmt_860/merge_stmt_1479_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_860/merge_stmt_1479_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_860/merge_stmt_1479_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_860/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_860/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_860/assign_stmt_1477/WPIPE_Block0_complete_1475_Update/$exit
      -- 
    ack_3846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1475_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(88)); -- 
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	16 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_req
      -- CP-element group 89: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1033_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1029/$exit
      -- 
    phi_stmt_1029_req_3857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1029_req_3857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(89), ack => phi_stmt_1029_req_0); -- 
    -- Element group zeropad3D_A_CP_2698_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2698_elements(16), ack => zeropad3D_A_CP_2698_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	16 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1036/$exit
      -- CP-element group 90: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1040_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_req
      -- 
    phi_stmt_1036_req_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1036_req_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(90), ack => phi_stmt_1036_req_0); -- 
    -- Element group zeropad3D_A_CP_2698_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2698_elements(16), ack => zeropad3D_A_CP_2698_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  transition  output  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	16 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_req
      -- CP-element group 91: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1047_konst_delay_trans
      -- CP-element group 91: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/phi_stmt_1043/$exit
      -- 
    phi_stmt_1043_req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1043_req_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(91), ack => phi_stmt_1043_req_0); -- 
    -- Element group zeropad3D_A_CP_2698_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2698_elements(16), ack => zeropad3D_A_CP_2698_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  join  transition  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	89 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	103 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_860/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(89) & zeropad3D_A_CP_2698_elements(90) & zeropad3D_A_CP_2698_elements(91);
      gj_zeropad3D_A_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Sample/$exit
      -- 
    ra_3893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/Update/$exit
      -- 
    ca_3898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	102 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_req
      -- CP-element group 95: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/type_cast_1035/$exit
      -- CP-element group 95: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/phi_stmt_1029_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1029/$exit
      -- 
    phi_stmt_1029_req_3899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1029_req_3899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(95), ack => phi_stmt_1029_req_1); -- 
    zeropad3D_A_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(93) & zeropad3D_A_CP_2698_elements(94);
      gj_zeropad3D_A_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/$exit
      -- 
    ra_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1042_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	1 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/ca
      -- CP-element group 97: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/$exit
      -- 
    ca_3921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1042_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_req
      -- CP-element group 98: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/$exit
      -- CP-element group 98: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/$exit
      -- CP-element group 98: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$exit
      -- CP-element group 98: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1036/$exit
      -- 
    phi_stmt_1036_req_3922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1036_req_3922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(98), ack => phi_stmt_1036_req_1); -- 
    zeropad3D_A_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(96) & zeropad3D_A_CP_2698_elements(97);
      gj_zeropad3D_A_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/ra
      -- 
    ra_3939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/ca
      -- 
    ca_3944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/$exit
      -- CP-element group 101: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/$exit
      -- CP-element group 101: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/phi_stmt_1043/phi_stmt_1043_req
      -- 
    phi_stmt_1043_req_3945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1043_req_3945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(101), ack => phi_stmt_1043_req_1); -- 
    zeropad3D_A_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(99) & zeropad3D_A_CP_2698_elements(100);
      gj_zeropad3D_A_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	95 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_860/ifx_xend170_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(95) & zeropad3D_A_CP_2698_elements(98) & zeropad3D_A_CP_2698_elements(101);
      gj_zeropad3D_A_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  merge  fork  transition  place  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	92 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	105 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_860/merge_stmt_1028_PhiReqMerge
      -- CP-element group 103: 	 branch_block_stmt_860/merge_stmt_1028_PhiAck/$entry
      -- 
    zeropad3D_A_CP_2698_elements(103) <= OrReduce(zeropad3D_A_CP_2698_elements(92) & zeropad3D_A_CP_2698_elements(102));
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_860/merge_stmt_1028_PhiAck/phi_stmt_1029_ack
      -- 
    phi_stmt_1029_ack_3950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1029_ack_0, ack => zeropad3D_A_CP_2698_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_860/merge_stmt_1028_PhiAck/phi_stmt_1036_ack
      -- 
    phi_stmt_1036_ack_3951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1036_ack_0, ack => zeropad3D_A_CP_2698_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_860/merge_stmt_1028_PhiAck/phi_stmt_1043_ack
      -- 
    phi_stmt_1043_ack_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1043_ack_0, ack => zeropad3D_A_CP_2698_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  place  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	18 
    -- CP-element group 107: 	17 
    -- CP-element group 107:  members (10) 
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/$entry
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062/type_cast_1054_update_start_
      -- CP-element group 107: 	 branch_block_stmt_860/merge_stmt_1028_PhiAck/$exit
      -- CP-element group 107: 	 branch_block_stmt_860/merge_stmt_1028__exit__
      -- CP-element group 107: 	 branch_block_stmt_860/assign_stmt_1055_to_assign_stmt_1062__entry__
      -- 
    cr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(107), ack => type_cast_1054_inst_req_1); -- 
    rr_3043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(107), ack => type_cast_1054_inst_req_0); -- 
    zeropad3D_A_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(104) & zeropad3D_A_CP_2698_elements(105) & zeropad3D_A_CP_2698_elements(106);
      gj_zeropad3D_A_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  merge  fork  transition  place  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	34 
    -- CP-element group 108: 	19 
    -- CP-element group 108: 	25 
    -- CP-element group 108: 	28 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	35 
    -- CP-element group 108: 	36 
    -- CP-element group 108: 	37 
    -- CP-element group 108: 	38 
    -- CP-element group 108: 	41 
    -- CP-element group 108: 	43 
    -- CP-element group 108: 	45 
    -- CP-element group 108: 	47 
    -- CP-element group 108:  members (33) 
      -- CP-element group 108: 	 branch_block_stmt_860/merge_stmt_1158_PhiReqMerge
      -- CP-element group 108: 	 branch_block_stmt_860/merge_stmt_1158__exit__
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214__entry__
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_update_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1162_Update/cr
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_update_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1167_Update/cr
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_update_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/type_cast_1201_Update/cr
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_update_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_update_start
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/array_obj_ref_1207_final_index_sum_regn_Update/req
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_complete/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/addr_of_1208_complete/req
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_update_start_
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/word_access_complete/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/word_access_complete/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_860/assign_stmt_1163_to_assign_stmt_1214/ptr_deref_1211_Update/word_access_complete/word_0/cr
      -- CP-element group 108: 	 branch_block_stmt_860/merge_stmt_1158_PhiAck/dummy
      -- CP-element group 108: 	 branch_block_stmt_860/merge_stmt_1158_PhiAck/$exit
      -- CP-element group 108: 	 branch_block_stmt_860/merge_stmt_1158_PhiAck/$entry
      -- 
    rr_3259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => type_cast_1162_inst_req_0); -- 
    cr_3264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => type_cast_1162_inst_req_1); -- 
    rr_3273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => type_cast_1167_inst_req_0); -- 
    cr_3278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => type_cast_1167_inst_req_1); -- 
    cr_3292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => type_cast_1201_inst_req_1); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => array_obj_ref_1207_index_offset_req_1); -- 
    req_3338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => addr_of_1208_final_reg_req_1); -- 
    cr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(108), ack => ptr_deref_1211_store_0_req_1); -- 
    zeropad3D_A_CP_2698_elements(108) <= OrReduce(zeropad3D_A_CP_2698_elements(34) & zeropad3D_A_CP_2698_elements(19) & zeropad3D_A_CP_2698_elements(25) & zeropad3D_A_CP_2698_elements(28));
    -- CP-element group 109:  merge  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	48 
    -- CP-element group 109: 	68 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	69 
    -- CP-element group 109: 	70 
    -- CP-element group 109:  members (13) 
      -- CP-element group 109: 	 branch_block_stmt_860/merge_stmt_1323_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_860/merge_stmt_1323__exit__
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341__entry__
      -- CP-element group 109: 	 branch_block_stmt_860/merge_stmt_1323_PhiAck/dummy
      -- CP-element group 109: 	 branch_block_stmt_860/merge_stmt_1323_PhiAck/$exit
      -- CP-element group 109: 	 branch_block_stmt_860/merge_stmt_1323_PhiAck/$entry
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/$entry
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_update_start_
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_860/assign_stmt_1328_to_assign_stmt_1341/type_cast_1327_Update/cr
      -- 
    rr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(109), ack => type_cast_1327_inst_req_0); -- 
    cr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(109), ack => type_cast_1327_inst_req_1); -- 
    zeropad3D_A_CP_2698_elements(109) <= OrReduce(zeropad3D_A_CP_2698_elements(48) & zeropad3D_A_CP_2698_elements(68));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	86 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Sample/$exit
      -- 
    ra_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1457_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	86 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Update/ca
      -- CP-element group 111: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/Update/$exit
      -- 
    ca_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1457_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	117 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/$exit
      -- CP-element group 112: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/$exit
      -- CP-element group 112: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/$exit
      -- CP-element group 112: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_req
      -- CP-element group 112: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1457/SplitProtocol/$exit
      -- 
    phi_stmt_1452_req_4078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1452_req_4078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(112), ack => phi_stmt_1452_req_1); -- 
    zeropad3D_A_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(110) & zeropad3D_A_CP_2698_elements(111);
      gj_zeropad3D_A_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Sample/$exit
      -- 
    ra_4095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	86 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Update/ca
      -- CP-element group 114: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/Update/$exit
      -- 
    ca_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_req
      -- CP-element group 115: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1463/$exit
      -- CP-element group 115: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1458/$exit
      -- 
    phi_stmt_1458_req_4101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1458_req_4101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(115), ack => phi_stmt_1458_req_1); -- 
    zeropad3D_A_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(113) & zeropad3D_A_CP_2698_elements(114);
      gj_zeropad3D_A_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  output  delay-element  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_req
      -- CP-element group 116: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1470_konst_delay_trans
      -- CP-element group 116: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/phi_stmt_1464/$exit
      -- 
    phi_stmt_1464_req_4109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1464_req_4109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(116), ack => phi_stmt_1464_req_1); -- 
    -- Element group zeropad3D_A_CP_2698_elements(116) is a control-delay.
    cp_element_116_delay: control_delay_element  generic map(name => " 116_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2698_elements(86), ack => zeropad3D_A_CP_2698_elements(116), clk => clk, reset =>reset);
    -- CP-element group 117:  join  transition  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	112 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	128 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_860/ifx_xelse138_ifx_xend170_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(112) & zeropad3D_A_CP_2698_elements(115) & zeropad3D_A_CP_2698_elements(116);
      gj_zeropad3D_A_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	71 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Sample/ra
      -- 
    ra_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	71 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Update/ca
      -- CP-element group 119: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/Update/$exit
      -- 
    ca_4134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	127 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/$exit
      -- CP-element group 120: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/type_cast_1455/SplitProtocol/$exit
      -- CP-element group 120: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_req
      -- CP-element group 120: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/phi_stmt_1452_sources/$exit
      -- CP-element group 120: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1452/$exit
      -- 
    phi_stmt_1452_req_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1452_req_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(120), ack => phi_stmt_1452_req_0); -- 
    zeropad3D_A_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(118) & zeropad3D_A_CP_2698_elements(119);
      gj_zeropad3D_A_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	71 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Sample/ra
      -- 
    ra_4152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1461_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	71 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Update/ca
      -- CP-element group 122: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/Update/$exit
      -- 
    ca_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1461_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	127 
    -- CP-element group 123:  members (5) 
      -- CP-element group 123: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/SplitProtocol/$exit
      -- CP-element group 123: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/type_cast_1461/$exit
      -- CP-element group 123: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_sources/$exit
      -- CP-element group 123: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/phi_stmt_1458_req
      -- CP-element group 123: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1458/$exit
      -- 
    phi_stmt_1458_req_4158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1458_req_4158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(123), ack => phi_stmt_1458_req_0); -- 
    zeropad3D_A_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(121) & zeropad3D_A_CP_2698_elements(122);
      gj_zeropad3D_A_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	71 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/$exit
      -- 
    ra_4175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_0, ack => zeropad3D_A_CP_2698_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	71 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/ca
      -- CP-element group 125: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/$exit
      -- 
    ca_4180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_1, ack => zeropad3D_A_CP_2698_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_req
      -- CP-element group 126: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/$exit
      -- CP-element group 126: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/$exit
      -- CP-element group 126: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/phi_stmt_1464/$exit
      -- 
    phi_stmt_1464_req_4181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1464_req_4181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2698_elements(126), ack => phi_stmt_1464_req_0); -- 
    zeropad3D_A_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(124) & zeropad3D_A_CP_2698_elements(125);
      gj_zeropad3D_A_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	120 
    -- CP-element group 127: 	123 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_860/ifx_xthen133_ifx_xend170_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(120) & zeropad3D_A_CP_2698_elements(123) & zeropad3D_A_CP_2698_elements(126);
      gj_zeropad3D_A_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  merge  fork  transition  place  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	117 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: 	130 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_860/merge_stmt_1451_PhiAck/$entry
      -- CP-element group 128: 	 branch_block_stmt_860/merge_stmt_1451_PhiReqMerge
      -- 
    zeropad3D_A_CP_2698_elements(128) <= OrReduce(zeropad3D_A_CP_2698_elements(117) & zeropad3D_A_CP_2698_elements(127));
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	132 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_860/merge_stmt_1451_PhiAck/phi_stmt_1452_ack
      -- 
    phi_stmt_1452_ack_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1452_ack_0, ack => zeropad3D_A_CP_2698_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_860/merge_stmt_1451_PhiAck/phi_stmt_1458_ack
      -- 
    phi_stmt_1458_ack_4187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1458_ack_0, ack => zeropad3D_A_CP_2698_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	128 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_860/merge_stmt_1451_PhiAck/phi_stmt_1464_ack
      -- 
    phi_stmt_1464_ack_4188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1464_ack_0, ack => zeropad3D_A_CP_2698_elements(131)); -- 
    -- CP-element group 132:  join  transition  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	129 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	1 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_860/merge_stmt_1451_PhiAck/$exit
      -- 
    zeropad3D_A_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2698_elements(129) & zeropad3D_A_CP_2698_elements(130) & zeropad3D_A_CP_2698_elements(131);
      gj_zeropad3D_A_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2698_elements(132), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1024_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1195_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1278_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1303_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_929_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_944_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_959_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_983_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_998_wire : std_logic_vector(31 downto 0);
    signal LOAD_pad_866_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_866_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom118_1289_resized : std_logic_vector(13 downto 0);
    signal R_idxprom118_1289_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom123_1314_resized : std_logic_vector(13 downto 0);
    signal R_idxprom123_1314_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1206_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1206_scaled : std_logic_vector(13 downto 0);
    signal add109_1266 : std_logic_vector(31 downto 0);
    signal add115_1271 : std_logic_vector(31 downto 0);
    signal add128_1334 : std_logic_vector(31 downto 0);
    signal add136_1354 : std_logic_vector(15 downto 0);
    signal add146_1390 : std_logic_vector(31 downto 0);
    signal add161_1439 : std_logic_vector(31 downto 0);
    signal add61_1146 : std_logic_vector(31 downto 0);
    signal add72_1183 : std_logic_vector(31 downto 0);
    signal add78_1188 : std_logic_vector(31 downto 0);
    signal add90_1246 : std_logic_vector(31 downto 0);
    signal add99_1251 : std_logic_vector(31 downto 0);
    signal add_1092 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1207_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1290_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1290_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1290_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1290_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1290_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1290_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1315_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1315_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1315_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1315_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1315_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1315_root_address : std_logic_vector(13 downto 0);
    signal arrayidx119_1292 : std_logic_vector(31 downto 0);
    signal arrayidx124_1317 : std_logic_vector(31 downto 0);
    signal arrayidx_1209 : std_logic_vector(31 downto 0);
    signal call_863 : std_logic_vector(15 downto 0);
    signal cmp131_1341 : std_logic_vector(0 downto 0);
    signal cmp147_1395 : std_logic_vector(0 downto 0);
    signal cmp162_1444 : std_logic_vector(0 downto 0);
    signal cmp45_1097 : std_logic_vector(0 downto 0);
    signal cmp52_1116 : std_logic_vector(0 downto 0);
    signal cmp62_1151 : std_logic_vector(0 downto 0);
    signal cmp_1062 : std_logic_vector(0 downto 0);
    signal conv127_1328 : std_logic_vector(31 downto 0);
    signal conv130_1000 : std_logic_vector(31 downto 0);
    signal conv141_1367 : std_logic_vector(31 downto 0);
    signal conv155_1416 : std_logic_vector(31 downto 0);
    signal conv23_931 : std_logic_vector(31 downto 0);
    signal conv27_946 : std_logic_vector(31 downto 0);
    signal conv29_961 : std_logic_vector(31 downto 0);
    signal conv36_1055 : std_logic_vector(31 downto 0);
    signal conv38_970 : std_logic_vector(31 downto 0);
    signal conv49_1109 : std_logic_vector(31 downto 0);
    signal conv66_1163 : std_logic_vector(31 downto 0);
    signal conv70_1168 : std_logic_vector(31 downto 0);
    signal conv74_985 : std_logic_vector(31 downto 0);
    signal conv82_1221 : std_logic_vector(31 downto 0);
    signal conv92_1026 : std_logic_vector(31 downto 0);
    signal div143_1385 : std_logic_vector(31 downto 0);
    signal div157_1434 : std_logic_vector(31 downto 0);
    signal div58_1141 : std_logic_vector(31 downto 0);
    signal div_1087 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1077 : std_logic_vector(31 downto 0);
    signal iNsTr_15_1375 : std_logic_vector(31 downto 0);
    signal iNsTr_16_1424 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1131 : std_logic_vector(31 downto 0);
    signal iNsTr_2_875 : std_logic_vector(31 downto 0);
    signal iNsTr_3_887 : std_logic_vector(31 downto 0);
    signal iNsTr_4_899 : std_logic_vector(31 downto 0);
    signal iNsTr_5_911 : std_logic_vector(31 downto 0);
    signal idxprom118_1285 : std_logic_vector(63 downto 0);
    signal idxprom123_1310 : std_logic_vector(63 downto 0);
    signal idxprom_1202 : std_logic_vector(63 downto 0);
    signal inc152_1399 : std_logic_vector(15 downto 0);
    signal inc152x_xix_x2_1404 : std_logic_vector(15 downto 0);
    signal inc_1362 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1452 : std_logic_vector(15 downto 0);
    signal ix_x2_1029 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1458 : std_logic_vector(15 downto 0);
    signal jx_x1_1036 : std_logic_vector(15 downto 0);
    signal jx_x2_1411 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1464 : std_logic_vector(15 downto 0);
    signal kx_x1_1043 : std_logic_vector(15 downto 0);
    signal mul108_1256 : std_logic_vector(31 downto 0);
    signal mul114_1261 : std_logic_vector(31 downto 0);
    signal mul30_966 : std_logic_vector(31 downto 0);
    signal mul71_1173 : std_logic_vector(31 downto 0);
    signal mul77_1178 : std_logic_vector(31 downto 0);
    signal mul89_1231 : std_logic_vector(31 downto 0);
    signal mul98_1241 : std_logic_vector(31 downto 0);
    signal mul_1012 : std_logic_vector(31 downto 0);
    signal ptr_deref_1080_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1080_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1080_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1080_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1080_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1134_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1134_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1134_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1134_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1134_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1211_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1211_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1211_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1211_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1211_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1211_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1295_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1295_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1295_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1295_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1295_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1319_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1319_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1319_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1319_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1319_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1319_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1378_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1378_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1378_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1378_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1378_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1427_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1427_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1427_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1427_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1427_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_878_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_878_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_878_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_878_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_878_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_890_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_890_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_890_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_890_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_890_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_902_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_902_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_902_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_902_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_902_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_914_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_914_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_914_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_914_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_914_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext172_952 : std_logic_vector(31 downto 0);
    signal sext173_1017 : std_logic_vector(31 downto 0);
    signal sext179_937 : std_logic_vector(31 downto 0);
    signal sext180_976 : std_logic_vector(31 downto 0);
    signal sext181_991 : std_logic_vector(31 downto 0);
    signal sext_921 : std_logic_vector(31 downto 0);
    signal shl_1006 : std_logic_vector(31 downto 0);
    signal shr117_1280 : std_logic_vector(31 downto 0);
    signal shr122_1305 : std_logic_vector(31 downto 0);
    signal shr_1197 : std_logic_vector(31 downto 0);
    signal sub97_1236 : std_logic_vector(31 downto 0);
    signal sub_1226 : std_logic_vector(31 downto 0);
    signal tmp11_903 : std_logic_vector(31 downto 0);
    signal tmp120_1296 : std_logic_vector(63 downto 0);
    signal tmp142_1379 : std_logic_vector(31 downto 0);
    signal tmp14_915 : std_logic_vector(31 downto 0);
    signal tmp156_1428 : std_logic_vector(31 downto 0);
    signal tmp2_879 : std_logic_vector(31 downto 0);
    signal tmp42_1081 : std_logic_vector(31 downto 0);
    signal tmp57_1135 : std_logic_vector(31 downto 0);
    signal tmp5_891 : std_logic_vector(31 downto 0);
    signal tmp_867 : std_logic_vector(7 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1020_wire : std_logic_vector(31 downto 0);
    signal type_cast_1023_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1033_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1035_wire : std_logic_vector(15 downto 0);
    signal type_cast_1040_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1042_wire : std_logic_vector(15 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1049_wire : std_logic_vector(15 downto 0);
    signal type_cast_1053_wire : std_logic_vector(31 downto 0);
    signal type_cast_1058_wire : std_logic_vector(31 downto 0);
    signal type_cast_1060_wire : std_logic_vector(31 downto 0);
    signal type_cast_1085_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1107_wire : std_logic_vector(31 downto 0);
    signal type_cast_1112_wire : std_logic_vector(31 downto 0);
    signal type_cast_1114_wire : std_logic_vector(31 downto 0);
    signal type_cast_1139_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1161_wire : std_logic_vector(31 downto 0);
    signal type_cast_1166_wire : std_logic_vector(31 downto 0);
    signal type_cast_1191_wire : std_logic_vector(31 downto 0);
    signal type_cast_1194_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1200_wire : std_logic_vector(63 downto 0);
    signal type_cast_1213_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1219_wire : std_logic_vector(31 downto 0);
    signal type_cast_1274_wire : std_logic_vector(31 downto 0);
    signal type_cast_1277_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1283_wire : std_logic_vector(63 downto 0);
    signal type_cast_1299_wire : std_logic_vector(31 downto 0);
    signal type_cast_1302_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1308_wire : std_logic_vector(63 downto 0);
    signal type_cast_1326_wire : std_logic_vector(31 downto 0);
    signal type_cast_1332_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1337_wire : std_logic_vector(31 downto 0);
    signal type_cast_1339_wire : std_logic_vector(31 downto 0);
    signal type_cast_1352_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1360_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1365_wire : std_logic_vector(31 downto 0);
    signal type_cast_1383_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1408_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1414_wire : std_logic_vector(31 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1455_wire : std_logic_vector(15 downto 0);
    signal type_cast_1457_wire : std_logic_vector(15 downto 0);
    signal type_cast_1461_wire : std_logic_vector(15 downto 0);
    signal type_cast_1463_wire : std_logic_vector(15 downto 0);
    signal type_cast_1467_wire : std_logic_vector(15 downto 0);
    signal type_cast_1470_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_919_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_925_wire : std_logic_vector(31 downto 0);
    signal type_cast_928_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_935_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_940_wire : std_logic_vector(31 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_950_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_955_wire : std_logic_vector(31 downto 0);
    signal type_cast_958_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_974_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_979_wire : std_logic_vector(31 downto 0);
    signal type_cast_982_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_989_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_994_wire : std_logic_vector(31 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_pad_866_word_address_0 <= "0";
    array_obj_ref_1207_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1207_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1207_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1207_resized_base_address <= "00000000000000";
    array_obj_ref_1290_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1290_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1290_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1290_resized_base_address <= "00000000000000";
    array_obj_ref_1315_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1315_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1315_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1315_resized_base_address <= "00000000000000";
    iNsTr_10_1077 <= "00000000000000000000000000000011";
    iNsTr_15_1375 <= "00000000000000000000000000000100";
    iNsTr_16_1424 <= "00000000000000000000000000000011";
    iNsTr_18_1131 <= "00000000000000000000000000000100";
    iNsTr_2_875 <= "00000000000000000000000000000101";
    iNsTr_3_887 <= "00000000000000000000000000000100";
    iNsTr_4_899 <= "00000000000000000000000000000101";
    iNsTr_5_911 <= "00000000000000000000000000000100";
    ptr_deref_1080_word_offset_0 <= "0000000";
    ptr_deref_1134_word_offset_0 <= "0000000";
    ptr_deref_1211_word_offset_0 <= "00000000000000";
    ptr_deref_1295_word_offset_0 <= "00000000000000";
    ptr_deref_1319_word_offset_0 <= "00000000000000";
    ptr_deref_1378_word_offset_0 <= "0000000";
    ptr_deref_1427_word_offset_0 <= "0000000";
    ptr_deref_878_word_offset_0 <= "0000000";
    ptr_deref_890_word_offset_0 <= "0000000";
    ptr_deref_902_word_offset_0 <= "0000000";
    ptr_deref_914_word_offset_0 <= "0000000";
    type_cast_1004_wire_constant <= "00000000000000000000000000000001";
    type_cast_1010_wire_constant <= "00000000000000000000000000010000";
    type_cast_1023_wire_constant <= "00000000000000000000000000010000";
    type_cast_1033_wire_constant <= "0000000000000000";
    type_cast_1040_wire_constant <= "0000000000000000";
    type_cast_1047_wire_constant <= "0000000000000000";
    type_cast_1085_wire_constant <= "00000000000000000000000000000001";
    type_cast_1139_wire_constant <= "00000000000000000000000000000001";
    type_cast_1194_wire_constant <= "00000000000000000000000000000010";
    type_cast_1213_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1277_wire_constant <= "00000000000000000000000000000010";
    type_cast_1302_wire_constant <= "00000000000000000000000000000010";
    type_cast_1332_wire_constant <= "00000000000000000000000000000100";
    type_cast_1352_wire_constant <= "0000000000000100";
    type_cast_1360_wire_constant <= "0000000000000001";
    type_cast_1383_wire_constant <= "00000000000000000000000000000001";
    type_cast_1408_wire_constant <= "0000000000000000";
    type_cast_1432_wire_constant <= "00000000000000000000000000000001";
    type_cast_1470_wire_constant <= "0000000000000000";
    type_cast_919_wire_constant <= "00000000000000000000000000010000";
    type_cast_928_wire_constant <= "00000000000000000000000000010000";
    type_cast_935_wire_constant <= "00000000000000000000000000010000";
    type_cast_943_wire_constant <= "00000000000000000000000000010000";
    type_cast_950_wire_constant <= "00000000000000000000000000010000";
    type_cast_958_wire_constant <= "00000000000000000000000000010000";
    type_cast_974_wire_constant <= "00000000000000000000000000010000";
    type_cast_982_wire_constant <= "00000000000000000000000000010000";
    type_cast_989_wire_constant <= "00000000000000000000000000010000";
    type_cast_997_wire_constant <= "00000000000000000000000000010000";
    phi_stmt_1029: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1033_wire_constant & type_cast_1035_wire;
      req <= phi_stmt_1029_req_0 & phi_stmt_1029_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1029",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1029_ack_0,
          idata => idata,
          odata => ix_x2_1029,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1029
    phi_stmt_1036: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1040_wire_constant & type_cast_1042_wire;
      req <= phi_stmt_1036_req_0 & phi_stmt_1036_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1036",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1036_ack_0,
          idata => idata,
          odata => jx_x1_1036,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1036
    phi_stmt_1043: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1047_wire_constant & type_cast_1049_wire;
      req <= phi_stmt_1043_req_0 & phi_stmt_1043_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1043",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1043_ack_0,
          idata => idata,
          odata => kx_x1_1043,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1043
    phi_stmt_1452: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1455_wire & type_cast_1457_wire;
      req <= phi_stmt_1452_req_0 & phi_stmt_1452_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1452",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1452_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1452,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1452
    phi_stmt_1458: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1461_wire & type_cast_1463_wire;
      req <= phi_stmt_1458_req_0 & phi_stmt_1458_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1458",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1458_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1458,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1458
    phi_stmt_1464: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1467_wire & type_cast_1470_wire_constant;
      req <= phi_stmt_1464_req_0 & phi_stmt_1464_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1464",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1464_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1464,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1464
    -- flow-through select operator MUX_1410_inst
    jx_x2_1411 <= type_cast_1408_wire_constant when (cmp147_1395(0) /=  '0') else inc_1362;
    addr_of_1208_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1208_final_reg_req_0;
      addr_of_1208_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1208_final_reg_req_1;
      addr_of_1208_final_reg_ack_1<= rack(0);
      addr_of_1208_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1208_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1207_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1291_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1291_final_reg_req_0;
      addr_of_1291_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1291_final_reg_req_1;
      addr_of_1291_final_reg_ack_1<= rack(0);
      addr_of_1291_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1291_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1290_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx119_1292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1316_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1316_final_reg_req_0;
      addr_of_1316_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1316_final_reg_req_1;
      addr_of_1316_final_reg_ack_1<= rack(0);
      addr_of_1316_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1316_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1315_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx124_1317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1020_inst
    process(sext173_1017) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext173_1017(31 downto 0);
      type_cast_1020_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1025_inst
    process(ASHR_i32_i32_1024_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1024_wire(31 downto 0);
      conv92_1026 <= tmp_var; -- 
    end process;
    type_cast_1035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1035_inst_req_0;
      type_cast_1035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1035_inst_req_1;
      type_cast_1035_inst_ack_1<= rack(0);
      type_cast_1035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1035_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1042_inst_req_0;
      type_cast_1042_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1042_inst_req_1;
      type_cast_1042_inst_ack_1<= rack(0);
      type_cast_1042_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1042_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1042_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1049_inst_req_0;
      type_cast_1049_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1049_inst_req_1;
      type_cast_1049_inst_ack_1<= rack(0);
      type_cast_1049_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1049_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1049_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1054_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1054_inst_req_0;
      type_cast_1054_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1054_inst_req_1;
      type_cast_1054_inst_ack_1<= rack(0);
      type_cast_1054_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1054_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1053_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_1055,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1058_inst
    process(conv36_1055) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_1055(31 downto 0);
      type_cast_1058_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1060_inst
    process(conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv38_970(31 downto 0);
      type_cast_1060_wire <= tmp_var; -- 
    end process;
    type_cast_1108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1108_inst_req_0;
      type_cast_1108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1108_inst_req_1;
      type_cast_1108_inst_ack_1<= rack(0);
      type_cast_1108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1107_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1112_inst
    process(conv49_1109) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_1109(31 downto 0);
      type_cast_1112_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1114_inst
    process(conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv38_970(31 downto 0);
      type_cast_1114_wire <= tmp_var; -- 
    end process;
    type_cast_1162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1162_inst_req_0;
      type_cast_1162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1162_inst_req_1;
      type_cast_1162_inst_ack_1<= rack(0);
      type_cast_1162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1161_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1166_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1191_inst
    process(add78_1188) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add78_1188(31 downto 0);
      type_cast_1191_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1196_inst
    process(ASHR_i32_i32_1195_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1195_wire(31 downto 0);
      shr_1197 <= tmp_var; -- 
    end process;
    type_cast_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1201_inst_req_0;
      type_cast_1201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1201_inst_req_1;
      type_cast_1201_inst_ack_1<= rack(0);
      type_cast_1201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1200_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1220_inst_req_0;
      type_cast_1220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1220_inst_req_1;
      type_cast_1220_inst_ack_1<= rack(0);
      type_cast_1220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1219_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1274_inst
    process(add99_1251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add99_1251(31 downto 0);
      type_cast_1274_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1279_inst
    process(ASHR_i32_i32_1278_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1278_wire(31 downto 0);
      shr117_1280 <= tmp_var; -- 
    end process;
    type_cast_1284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1284_inst_req_0;
      type_cast_1284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1284_inst_req_1;
      type_cast_1284_inst_ack_1<= rack(0);
      type_cast_1284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1283_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom118_1285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1299_inst
    process(add115_1271) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add115_1271(31 downto 0);
      type_cast_1299_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1304_inst
    process(ASHR_i32_i32_1303_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1303_wire(31 downto 0);
      shr122_1305 <= tmp_var; -- 
    end process;
    type_cast_1309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1309_inst_req_0;
      type_cast_1309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1309_inst_req_1;
      type_cast_1309_inst_ack_1<= rack(0);
      type_cast_1309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1308_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom123_1310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1327_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1327_inst_req_0;
      type_cast_1327_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1327_inst_req_1;
      type_cast_1327_inst_ack_1<= rack(0);
      type_cast_1327_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1327_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1326_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_1328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1337_inst
    process(add128_1334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add128_1334(31 downto 0);
      type_cast_1337_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1339_inst
    process(conv130_1000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv130_1000(31 downto 0);
      type_cast_1339_wire <= tmp_var; -- 
    end process;
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1365_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_1367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1398_inst_req_0;
      type_cast_1398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1398_inst_req_1;
      type_cast_1398_inst_ack_1<= rack(0);
      type_cast_1398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp147_1395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc152_1399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1415_inst_req_0;
      type_cast_1415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1415_inst_req_1;
      type_cast_1415_inst_ack_1<= rack(0);
      type_cast_1415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1414_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_1416,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1455_inst_req_0;
      type_cast_1455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1455_inst_req_1;
      type_cast_1455_inst_ack_1<= rack(0);
      type_cast_1455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1455_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1457_inst_req_0;
      type_cast_1457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1457_inst_req_1;
      type_cast_1457_inst_ack_1<= rack(0);
      type_cast_1457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc152x_xix_x2_1404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1457_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1461_inst_req_0;
      type_cast_1461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1461_inst_req_1;
      type_cast_1461_inst_ack_1<= rack(0);
      type_cast_1461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_1036,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1461_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1463_inst_req_0;
      type_cast_1463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1463_inst_req_1;
      type_cast_1463_inst_ack_1<= rack(0);
      type_cast_1463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1463_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1411,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1463_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1467_inst_req_0;
      type_cast_1467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1467_inst_req_1;
      type_cast_1467_inst_ack_1<= rack(0);
      type_cast_1467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add136_1354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1467_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_925_inst
    process(sext_921) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_921(31 downto 0);
      type_cast_925_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_930_inst
    process(ASHR_i32_i32_929_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_929_wire(31 downto 0);
      conv23_931 <= tmp_var; -- 
    end process;
    -- interlock type_cast_940_inst
    process(sext179_937) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext179_937(31 downto 0);
      type_cast_940_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_945_inst
    process(ASHR_i32_i32_944_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_944_wire(31 downto 0);
      conv27_946 <= tmp_var; -- 
    end process;
    -- interlock type_cast_955_inst
    process(sext172_952) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext172_952(31 downto 0);
      type_cast_955_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_960_inst
    process(ASHR_i32_i32_959_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_959_wire(31 downto 0);
      conv29_961 <= tmp_var; -- 
    end process;
    type_cast_969_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_969_inst_req_0;
      type_cast_969_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_969_inst_req_1;
      type_cast_969_inst_ack_1<= rack(0);
      type_cast_969_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_969_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_970,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_979_inst
    process(sext180_976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext180_976(31 downto 0);
      type_cast_979_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_984_inst
    process(ASHR_i32_i32_983_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_983_wire(31 downto 0);
      conv74_985 <= tmp_var; -- 
    end process;
    -- interlock type_cast_994_inst
    process(sext181_991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext181_991(31 downto 0);
      type_cast_994_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_999_inst
    process(ASHR_i32_i32_998_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_998_wire(31 downto 0);
      conv130_1000 <= tmp_var; -- 
    end process;
    -- equivalence LOAD_pad_866_gather_scatter
    process(LOAD_pad_866_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_866_data_0;
      ov(7 downto 0) := iv;
      tmp_867 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1207_index_1_rename
    process(R_idxprom_1206_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1206_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1206_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1207_index_1_resize
    process(idxprom_1202) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1202;
      ov := iv(13 downto 0);
      R_idxprom_1206_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1207_root_address_inst
    process(array_obj_ref_1207_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1207_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1207_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1290_index_1_rename
    process(R_idxprom118_1289_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom118_1289_resized;
      ov(13 downto 0) := iv;
      R_idxprom118_1289_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1290_index_1_resize
    process(idxprom118_1285) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom118_1285;
      ov := iv(13 downto 0);
      R_idxprom118_1289_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1290_root_address_inst
    process(array_obj_ref_1290_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1290_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1290_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1315_index_1_rename
    process(R_idxprom123_1314_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom123_1314_resized;
      ov(13 downto 0) := iv;
      R_idxprom123_1314_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1315_index_1_resize
    process(idxprom123_1310) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom123_1310;
      ov := iv(13 downto 0);
      R_idxprom123_1314_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1315_root_address_inst
    process(array_obj_ref_1315_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1315_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1315_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1080_addr_0
    process(ptr_deref_1080_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1080_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1080_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1080_base_resize
    process(iNsTr_10_1077) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1077;
      ov := iv(6 downto 0);
      ptr_deref_1080_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1080_gather_scatter
    process(ptr_deref_1080_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1080_data_0;
      ov(31 downto 0) := iv;
      tmp42_1081 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1080_root_address_inst
    process(ptr_deref_1080_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1080_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1080_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1134_addr_0
    process(ptr_deref_1134_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1134_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1134_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1134_base_resize
    process(iNsTr_18_1131) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_1131;
      ov := iv(6 downto 0);
      ptr_deref_1134_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1134_gather_scatter
    process(ptr_deref_1134_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1134_data_0;
      ov(31 downto 0) := iv;
      tmp57_1135 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1134_root_address_inst
    process(ptr_deref_1134_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1134_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1134_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1211_addr_0
    process(ptr_deref_1211_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1211_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1211_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1211_base_resize
    process(arrayidx_1209) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1209;
      ov := iv(13 downto 0);
      ptr_deref_1211_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1211_gather_scatter
    process(type_cast_1213_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1213_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1211_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1211_root_address_inst
    process(ptr_deref_1211_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1211_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1211_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1295_addr_0
    process(ptr_deref_1295_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1295_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1295_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1295_base_resize
    process(arrayidx119_1292) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx119_1292;
      ov := iv(13 downto 0);
      ptr_deref_1295_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1295_gather_scatter
    process(ptr_deref_1295_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1295_data_0;
      ov(63 downto 0) := iv;
      tmp120_1296 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1295_root_address_inst
    process(ptr_deref_1295_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1295_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1295_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1319_addr_0
    process(ptr_deref_1319_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1319_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1319_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1319_base_resize
    process(arrayidx124_1317) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx124_1317;
      ov := iv(13 downto 0);
      ptr_deref_1319_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1319_gather_scatter
    process(tmp120_1296) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp120_1296;
      ov(63 downto 0) := iv;
      ptr_deref_1319_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1319_root_address_inst
    process(ptr_deref_1319_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1319_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1319_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1378_addr_0
    process(ptr_deref_1378_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1378_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1378_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1378_base_resize
    process(iNsTr_15_1375) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_1375;
      ov := iv(6 downto 0);
      ptr_deref_1378_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1378_gather_scatter
    process(ptr_deref_1378_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1378_data_0;
      ov(31 downto 0) := iv;
      tmp142_1379 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1378_root_address_inst
    process(ptr_deref_1378_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1378_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1378_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1427_addr_0
    process(ptr_deref_1427_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1427_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1427_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1427_base_resize
    process(iNsTr_16_1424) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_16_1424;
      ov := iv(6 downto 0);
      ptr_deref_1427_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1427_gather_scatter
    process(ptr_deref_1427_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1427_data_0;
      ov(31 downto 0) := iv;
      tmp156_1428 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1427_root_address_inst
    process(ptr_deref_1427_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1427_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1427_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_878_addr_0
    process(ptr_deref_878_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_878_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_878_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_878_base_resize
    process(iNsTr_2_875) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_875;
      ov := iv(6 downto 0);
      ptr_deref_878_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_878_gather_scatter
    process(ptr_deref_878_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_878_data_0;
      ov(31 downto 0) := iv;
      tmp2_879 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_878_root_address_inst
    process(ptr_deref_878_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_878_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_878_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_890_addr_0
    process(ptr_deref_890_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_890_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_890_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_890_base_resize
    process(iNsTr_3_887) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_887;
      ov := iv(6 downto 0);
      ptr_deref_890_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_890_gather_scatter
    process(ptr_deref_890_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_890_data_0;
      ov(31 downto 0) := iv;
      tmp5_891 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_890_root_address_inst
    process(ptr_deref_890_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_890_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_890_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_902_addr_0
    process(ptr_deref_902_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_902_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_902_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_902_base_resize
    process(iNsTr_4_899) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_899;
      ov := iv(6 downto 0);
      ptr_deref_902_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_902_gather_scatter
    process(ptr_deref_902_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_902_data_0;
      ov(31 downto 0) := iv;
      tmp11_903 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_902_root_address_inst
    process(ptr_deref_902_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_902_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_902_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_914_addr_0
    process(ptr_deref_914_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_914_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_914_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_914_base_resize
    process(iNsTr_5_911) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_911;
      ov := iv(6 downto 0);
      ptr_deref_914_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_914_gather_scatter
    process(ptr_deref_914_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_914_data_0;
      ov(31 downto 0) := iv;
      tmp14_915 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_914_root_address_inst
    process(ptr_deref_914_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_914_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_914_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1063_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1062;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1063_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1063_branch_req_0,
          ack0 => if_stmt_1063_branch_ack_0,
          ack1 => if_stmt_1063_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1098_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp45_1097;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1098_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1098_branch_req_0,
          ack0 => if_stmt_1098_branch_ack_0,
          ack1 => if_stmt_1098_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1117_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp52_1116;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1117_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1117_branch_req_0,
          ack0 => if_stmt_1117_branch_ack_0,
          ack1 => if_stmt_1117_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1152_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp62_1151;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1152_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1152_branch_req_0,
          ack0 => if_stmt_1152_branch_ack_0,
          ack1 => if_stmt_1152_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1342_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp131_1341;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1342_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1342_branch_req_0,
          ack0 => if_stmt_1342_branch_ack_0,
          ack1 => if_stmt_1342_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1445_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp162_1444;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1445_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1445_branch_req_0,
          ack0 => if_stmt_1445_branch_ack_0,
          ack1 => if_stmt_1445_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1353_inst
    process(kx_x1_1043) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_1043, type_cast_1352_wire_constant, tmp_var);
      add136_1354 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1361_inst
    process(jx_x1_1036) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_1036, type_cast_1360_wire_constant, tmp_var);
      inc_1362 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1403_inst
    process(inc152_1399, ix_x2_1029) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc152_1399, ix_x2_1029, tmp_var);
      inc152x_xix_x2_1404 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1091_inst
    process(div_1087, conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div_1087, conv38_970, tmp_var);
      add_1092 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1145_inst
    process(div58_1141, conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div58_1141, conv38_970, tmp_var);
      add61_1146 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1182_inst
    process(mul71_1173, mul77_1178) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul71_1173, mul77_1178, tmp_var);
      add72_1183 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1187_inst
    process(add72_1183, conv66_1163) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add72_1183, conv66_1163, tmp_var);
      add78_1188 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1245_inst
    process(conv82_1221, mul98_1241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv82_1221, mul98_1241, tmp_var);
      add90_1246 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1250_inst
    process(add90_1246, mul89_1231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add90_1246, mul89_1231, tmp_var);
      add99_1251 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1265_inst
    process(mul108_1256, mul114_1261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul108_1256, mul114_1261, tmp_var);
      add109_1266 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1270_inst
    process(add109_1266, conv82_1221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add109_1266, conv82_1221, tmp_var);
      add115_1271 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1333_inst
    process(conv127_1328) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv127_1328, type_cast_1332_wire_constant, tmp_var);
      add128_1334 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1389_inst
    process(div143_1385, shl_1006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div143_1385, shl_1006, tmp_var);
      add146_1390 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1438_inst
    process(div157_1434, shl_1006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div157_1434, shl_1006, tmp_var);
      add161_1439 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1024_inst
    process(type_cast_1020_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1020_wire, type_cast_1023_wire_constant, tmp_var);
      ASHR_i32_i32_1024_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1195_inst
    process(type_cast_1191_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1191_wire, type_cast_1194_wire_constant, tmp_var);
      ASHR_i32_i32_1195_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1278_inst
    process(type_cast_1274_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1274_wire, type_cast_1277_wire_constant, tmp_var);
      ASHR_i32_i32_1278_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1303_inst
    process(type_cast_1299_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1299_wire, type_cast_1302_wire_constant, tmp_var);
      ASHR_i32_i32_1303_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_929_inst
    process(type_cast_925_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_925_wire, type_cast_928_wire_constant, tmp_var);
      ASHR_i32_i32_929_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_944_inst
    process(type_cast_940_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_940_wire, type_cast_943_wire_constant, tmp_var);
      ASHR_i32_i32_944_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_959_inst
    process(type_cast_955_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_955_wire, type_cast_958_wire_constant, tmp_var);
      ASHR_i32_i32_959_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_983_inst
    process(type_cast_979_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_979_wire, type_cast_982_wire_constant, tmp_var);
      ASHR_i32_i32_983_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_998_inst
    process(type_cast_994_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_994_wire, type_cast_997_wire_constant, tmp_var);
      ASHR_i32_i32_998_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1394_inst
    process(conv141_1367, add146_1390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv141_1367, add146_1390, tmp_var);
      cmp147_1395 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1443_inst
    process(conv155_1416, add161_1439) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv155_1416, add161_1439, tmp_var);
      cmp162_1444 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1086_inst
    process(tmp42_1081) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp42_1081, type_cast_1085_wire_constant, tmp_var);
      div_1087 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1140_inst
    process(tmp57_1135) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp57_1135, type_cast_1139_wire_constant, tmp_var);
      div58_1141 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1384_inst
    process(tmp142_1379) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp142_1379, type_cast_1383_wire_constant, tmp_var);
      div143_1385 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1433_inst
    process(tmp156_1428) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp156_1428, type_cast_1432_wire_constant, tmp_var);
      div157_1434 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1016_inst
    process(mul_1012, conv23_931) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1012, conv23_931, tmp_var);
      sext173_1017 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1172_inst
    process(conv70_1168, conv27_946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv70_1168, conv27_946, tmp_var);
      mul71_1173 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1177_inst
    process(conv36_1055, conv74_985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv36_1055, conv74_985, tmp_var);
      mul77_1178 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1230_inst
    process(sub_1226, conv130_1000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1226, conv130_1000, tmp_var);
      mul89_1231 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1240_inst
    process(sub97_1236, conv92_1026) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub97_1236, conv92_1026, tmp_var);
      mul98_1241 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1255_inst
    process(conv49_1109, conv27_946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv49_1109, conv27_946, tmp_var);
      mul108_1256 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1260_inst
    process(conv36_1055, conv74_985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv36_1055, conv74_985, tmp_var);
      mul114_1261 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_965_inst
    process(conv29_961, conv27_946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv29_961, conv27_946, tmp_var);
      mul30_966 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1005_inst
    process(conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv38_970, type_cast_1004_wire_constant, tmp_var);
      shl_1006 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1011_inst
    process(tmp2_879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp2_879, type_cast_1010_wire_constant, tmp_var);
      mul_1012 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_920_inst
    process(tmp5_891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp5_891, type_cast_919_wire_constant, tmp_var);
      sext_921 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_936_inst
    process(tmp11_903) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp11_903, type_cast_935_wire_constant, tmp_var);
      sext179_937 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_951_inst
    process(tmp14_915) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp14_915, type_cast_950_wire_constant, tmp_var);
      sext172_952 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_975_inst
    process(mul30_966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul30_966, type_cast_974_wire_constant, tmp_var);
      sext180_976 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_990_inst
    process(tmp2_879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp2_879, type_cast_989_wire_constant, tmp_var);
      sext181_991 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1061_inst
    process(type_cast_1058_wire, type_cast_1060_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1058_wire, type_cast_1060_wire, tmp_var);
      cmp_1062 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1115_inst
    process(type_cast_1112_wire, type_cast_1114_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1112_wire, type_cast_1114_wire, tmp_var);
      cmp52_1116 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1340_inst
    process(type_cast_1337_wire, type_cast_1339_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1337_wire, type_cast_1339_wire, tmp_var);
      cmp131_1341 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1225_inst
    process(conv49_1109, conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv49_1109, conv38_970, tmp_var);
      sub_1226 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1235_inst
    process(conv36_1055, conv38_970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv36_1055, conv38_970, tmp_var);
      sub97_1236 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1096_inst
    process(conv36_1055, add_1092) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv36_1055, add_1092, tmp_var);
      cmp45_1097 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1150_inst
    process(conv49_1109, add61_1146) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv49_1109, add61_1146, tmp_var);
      cmp62_1151 <= tmp_var; --
    end process;
    -- shared split operator group (51) : array_obj_ref_1207_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1206_scaled;
      array_obj_ref_1207_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1207_index_offset_req_0;
      array_obj_ref_1207_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1207_index_offset_req_1;
      array_obj_ref_1207_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : array_obj_ref_1290_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom118_1289_scaled;
      array_obj_ref_1290_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1290_index_offset_req_0;
      array_obj_ref_1290_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1290_index_offset_req_1;
      array_obj_ref_1290_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : array_obj_ref_1315_index_offset 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom123_1314_scaled;
      array_obj_ref_1315_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1315_index_offset_req_0;
      array_obj_ref_1315_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1315_index_offset_req_1;
      array_obj_ref_1315_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- unary operator type_cast_1053_inst
    process(ix_x2_1029) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_1029, tmp_var);
      type_cast_1053_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1107_inst
    process(jx_x1_1036) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1036, tmp_var);
      type_cast_1107_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1161_inst
    process(kx_x1_1043) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1043, tmp_var);
      type_cast_1161_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1166_inst
    process(jx_x1_1036) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1036, tmp_var);
      type_cast_1166_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1200_inst
    process(shr_1197) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1197, tmp_var);
      type_cast_1200_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1219_inst
    process(kx_x1_1043) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1043, tmp_var);
      type_cast_1219_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1283_inst
    process(shr117_1280) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr117_1280, tmp_var);
      type_cast_1283_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1308_inst
    process(shr122_1305) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr122_1305, tmp_var);
      type_cast_1308_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1326_inst
    process(kx_x1_1043) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1043, tmp_var);
      type_cast_1326_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1365_inst
    process(inc_1362) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1362, tmp_var);
      type_cast_1365_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1414_inst
    process(inc152x_xix_x2_1404) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc152x_xix_x2_1404, tmp_var);
      type_cast_1414_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_pad_866_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_pad_866_load_0_req_0;
      LOAD_pad_866_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_pad_866_load_0_req_1;
      LOAD_pad_866_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_866_word_address_0;
      LOAD_pad_866_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(0 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1378_load_0 ptr_deref_1427_load_0 ptr_deref_878_load_0 ptr_deref_890_load_0 ptr_deref_1080_load_0 ptr_deref_1134_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(41 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_1378_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1427_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_878_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_890_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1080_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1134_load_0_req_0;
      ptr_deref_1378_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1427_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_878_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_890_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1080_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1134_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_1378_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1427_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_878_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_890_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1080_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1134_load_0_req_1;
      ptr_deref_1378_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1427_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_878_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_890_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1080_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1134_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1378_word_address_0 & ptr_deref_1427_word_address_0 & ptr_deref_878_word_address_0 & ptr_deref_890_word_address_0 & ptr_deref_1080_word_address_0 & ptr_deref_1134_word_address_0;
      ptr_deref_1378_data_0 <= data_out(191 downto 160);
      ptr_deref_1427_data_0 <= data_out(159 downto 128);
      ptr_deref_878_data_0 <= data_out(127 downto 96);
      ptr_deref_890_data_0 <= data_out(95 downto 64);
      ptr_deref_1080_data_0 <= data_out(63 downto 32);
      ptr_deref_1134_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1295_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1295_load_0_req_0;
      ptr_deref_1295_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1295_load_0_req_1;
      ptr_deref_1295_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1295_word_address_0;
      ptr_deref_1295_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_902_load_0 ptr_deref_914_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_902_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_914_load_0_req_0;
      ptr_deref_902_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_914_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_902_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_914_load_0_req_1;
      ptr_deref_902_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_914_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_902_word_address_0 & ptr_deref_914_word_address_0;
      ptr_deref_902_data_0 <= data_out(63 downto 32);
      ptr_deref_914_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(6 downto 0),
          mtag => memory_space_4_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_1211_store_0 ptr_deref_1319_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1211_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1319_store_0_req_0;
      ptr_deref_1211_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1319_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1211_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1319_store_0_req_1;
      ptr_deref_1211_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1319_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1211_word_address_0 & ptr_deref_1319_word_address_0;
      data_in <= ptr_deref_1211_data_0 & ptr_deref_1319_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_starting_862_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_starting_862_inst_req_0;
      RPIPE_Block0_starting_862_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_starting_862_inst_req_1;
      RPIPE_Block0_starting_862_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_863 <= data_out(15 downto 0);
      Block0_starting_read_0_gI: SplitGuardInterface generic map(name => "Block0_starting_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block0_starting_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_starting_pipe_read_req(0),
          oack => Block0_starting_pipe_read_ack(0),
          odata => Block0_starting_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_complete_1475_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_complete_1475_inst_req_0;
      WPIPE_Block0_complete_1475_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_complete_1475_inst_req_1;
      WPIPE_Block0_complete_1475_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_863;
      Block0_complete_write_0_gI: SplitGuardInterface generic map(name => "Block0_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_complete", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_complete_pipe_write_req(0),
          oack => Block0_complete_pipe_write_ack(0),
          odata => Block0_complete_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_A_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_B is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block1_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_B;
architecture zeropad3D_B_arch of zeropad3D_B is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_B_CP_4205_start: Boolean;
  signal zeropad3D_B_CP_4205_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_pad_1511_load_0_req_1 : boolean;
  signal LOAD_pad_1511_load_0_req_0 : boolean;
  signal ptr_deref_1523_load_0_req_0 : boolean;
  signal phi_stmt_1646_req_0 : boolean;
  signal ptr_deref_1523_load_0_ack_0 : boolean;
  signal ptr_deref_1523_load_0_req_1 : boolean;
  signal ptr_deref_1498_load_0_req_1 : boolean;
  signal ptr_deref_1498_load_0_ack_1 : boolean;
  signal type_cast_1508_inst_ack_1 : boolean;
  signal type_cast_1508_inst_ack_0 : boolean;
  signal LOAD_pad_1511_load_0_ack_1 : boolean;
  signal ptr_deref_1523_load_0_ack_1 : boolean;
  signal type_cast_1508_inst_req_1 : boolean;
  signal LOAD_pad_1511_load_0_ack_0 : boolean;
  signal RPIPE_Block1_starting_1485_inst_req_0 : boolean;
  signal type_cast_1508_inst_req_0 : boolean;
  signal type_cast_1658_inst_ack_0 : boolean;
  signal ptr_deref_1547_load_0_req_1 : boolean;
  signal ptr_deref_1547_load_0_ack_1 : boolean;
  signal phi_stmt_2055_ack_0 : boolean;
  signal ptr_deref_1547_load_0_req_0 : boolean;
  signal ptr_deref_1547_load_0_ack_0 : boolean;
  signal phi_stmt_2067_req_1 : boolean;
  signal phi_stmt_2061_req_0 : boolean;
  signal ptr_deref_1535_load_0_req_1 : boolean;
  signal ptr_deref_1535_load_0_ack_1 : boolean;
  signal phi_stmt_2067_ack_0 : boolean;
  signal ptr_deref_1498_load_0_ack_0 : boolean;
  signal RPIPE_Block1_starting_1485_inst_ack_1 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal ptr_deref_1535_load_0_req_0 : boolean;
  signal ptr_deref_1498_load_0_req_0 : boolean;
  signal RPIPE_Block1_starting_1485_inst_req_1 : boolean;
  signal ptr_deref_1535_load_0_ack_0 : boolean;
  signal type_cast_1665_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1485_inst_ack_0 : boolean;
  signal phi_stmt_2055_req_1 : boolean;
  signal type_cast_2064_inst_ack_1 : boolean;
  signal type_cast_2060_inst_ack_1 : boolean;
  signal type_cast_1670_inst_req_0 : boolean;
  signal type_cast_1670_inst_ack_0 : boolean;
  signal type_cast_2060_inst_req_1 : boolean;
  signal type_cast_1670_inst_req_1 : boolean;
  signal phi_stmt_2061_req_1 : boolean;
  signal type_cast_1670_inst_ack_1 : boolean;
  signal phi_stmt_2061_ack_0 : boolean;
  signal if_stmt_1679_branch_req_0 : boolean;
  signal if_stmt_1679_branch_ack_1 : boolean;
  signal if_stmt_1679_branch_ack_0 : boolean;
  signal ptr_deref_1696_load_0_req_0 : boolean;
  signal ptr_deref_1696_load_0_ack_0 : boolean;
  signal ptr_deref_1696_load_0_req_1 : boolean;
  signal ptr_deref_1696_load_0_ack_1 : boolean;
  signal if_stmt_1714_branch_req_0 : boolean;
  signal if_stmt_1714_branch_ack_1 : boolean;
  signal if_stmt_1714_branch_ack_0 : boolean;
  signal type_cast_1724_inst_req_0 : boolean;
  signal type_cast_1724_inst_ack_0 : boolean;
  signal type_cast_1724_inst_req_1 : boolean;
  signal type_cast_1724_inst_ack_1 : boolean;
  signal if_stmt_1733_branch_req_0 : boolean;
  signal if_stmt_1733_branch_ack_1 : boolean;
  signal if_stmt_1733_branch_ack_0 : boolean;
  signal ptr_deref_1750_load_0_req_0 : boolean;
  signal ptr_deref_1750_load_0_ack_0 : boolean;
  signal ptr_deref_1750_load_0_req_1 : boolean;
  signal ptr_deref_1750_load_0_ack_1 : boolean;
  signal if_stmt_1762_branch_req_0 : boolean;
  signal if_stmt_1762_branch_ack_1 : boolean;
  signal if_stmt_1762_branch_ack_0 : boolean;
  signal type_cast_1772_inst_req_0 : boolean;
  signal type_cast_1772_inst_ack_0 : boolean;
  signal type_cast_1772_inst_req_1 : boolean;
  signal type_cast_1772_inst_ack_1 : boolean;
  signal type_cast_1777_inst_req_0 : boolean;
  signal type_cast_1777_inst_ack_0 : boolean;
  signal type_cast_1777_inst_req_1 : boolean;
  signal type_cast_1777_inst_ack_1 : boolean;
  signal type_cast_1811_inst_req_0 : boolean;
  signal type_cast_1811_inst_ack_0 : boolean;
  signal type_cast_1811_inst_req_1 : boolean;
  signal type_cast_1811_inst_ack_1 : boolean;
  signal type_cast_2064_inst_req_1 : boolean;
  signal phi_stmt_1653_req_0 : boolean;
  signal array_obj_ref_1817_index_offset_req_0 : boolean;
  signal type_cast_2066_inst_ack_1 : boolean;
  signal array_obj_ref_1817_index_offset_ack_0 : boolean;
  signal type_cast_2066_inst_req_1 : boolean;
  signal array_obj_ref_1817_index_offset_req_1 : boolean;
  signal array_obj_ref_1817_index_offset_ack_1 : boolean;
  signal type_cast_1665_inst_req_0 : boolean;
  signal addr_of_1818_final_reg_req_0 : boolean;
  signal addr_of_1818_final_reg_ack_0 : boolean;
  signal type_cast_2066_inst_ack_0 : boolean;
  signal addr_of_1818_final_reg_req_1 : boolean;
  signal addr_of_1818_final_reg_ack_1 : boolean;
  signal type_cast_2064_inst_ack_0 : boolean;
  signal type_cast_2064_inst_req_0 : boolean;
  signal type_cast_2066_inst_req_0 : boolean;
  signal type_cast_1658_inst_req_0 : boolean;
  signal ptr_deref_1821_store_0_req_0 : boolean;
  signal ptr_deref_1821_store_0_ack_0 : boolean;
  signal ptr_deref_1821_store_0_req_1 : boolean;
  signal ptr_deref_1821_store_0_ack_1 : boolean;
  signal type_cast_2060_inst_ack_0 : boolean;
  signal type_cast_1830_inst_req_0 : boolean;
  signal type_cast_1830_inst_ack_0 : boolean;
  signal type_cast_2060_inst_req_0 : boolean;
  signal type_cast_1830_inst_req_1 : boolean;
  signal type_cast_1830_inst_ack_1 : boolean;
  signal type_cast_1656_inst_ack_1 : boolean;
  signal type_cast_1894_inst_req_0 : boolean;
  signal type_cast_1894_inst_ack_0 : boolean;
  signal type_cast_1894_inst_req_1 : boolean;
  signal type_cast_1894_inst_ack_1 : boolean;
  signal phi_stmt_2055_req_0 : boolean;
  signal type_cast_2058_inst_ack_1 : boolean;
  signal type_cast_1656_inst_req_1 : boolean;
  signal array_obj_ref_1900_index_offset_req_0 : boolean;
  signal array_obj_ref_1900_index_offset_ack_0 : boolean;
  signal array_obj_ref_1900_index_offset_req_1 : boolean;
  signal array_obj_ref_1900_index_offset_ack_1 : boolean;
  signal addr_of_1901_final_reg_req_0 : boolean;
  signal addr_of_1901_final_reg_ack_0 : boolean;
  signal addr_of_1901_final_reg_req_1 : boolean;
  signal addr_of_1901_final_reg_ack_1 : boolean;
  signal type_cast_2058_inst_req_1 : boolean;
  signal type_cast_2058_inst_ack_0 : boolean;
  signal type_cast_2058_inst_req_0 : boolean;
  signal ptr_deref_1905_load_0_req_0 : boolean;
  signal ptr_deref_1905_load_0_ack_0 : boolean;
  signal ptr_deref_1905_load_0_req_1 : boolean;
  signal ptr_deref_1905_load_0_ack_1 : boolean;
  signal phi_stmt_2067_req_0 : boolean;
  signal type_cast_2070_inst_ack_1 : boolean;
  signal phi_stmt_1659_ack_0 : boolean;
  signal phi_stmt_1653_ack_0 : boolean;
  signal type_cast_2070_inst_req_1 : boolean;
  signal type_cast_1919_inst_req_0 : boolean;
  signal type_cast_1919_inst_ack_0 : boolean;
  signal type_cast_1656_inst_ack_0 : boolean;
  signal type_cast_1919_inst_req_1 : boolean;
  signal type_cast_1919_inst_ack_1 : boolean;
  signal phi_stmt_1659_req_1 : boolean;
  signal phi_stmt_1646_ack_0 : boolean;
  signal phi_stmt_1646_req_1 : boolean;
  signal type_cast_1652_inst_ack_1 : boolean;
  signal type_cast_1652_inst_req_1 : boolean;
  signal type_cast_1652_inst_ack_0 : boolean;
  signal type_cast_1656_inst_req_0 : boolean;
  signal type_cast_1652_inst_req_0 : boolean;
  signal array_obj_ref_1925_index_offset_req_0 : boolean;
  signal array_obj_ref_1925_index_offset_ack_0 : boolean;
  signal array_obj_ref_1925_index_offset_req_1 : boolean;
  signal array_obj_ref_1925_index_offset_ack_1 : boolean;
  signal type_cast_2070_inst_ack_0 : boolean;
  signal addr_of_1926_final_reg_req_0 : boolean;
  signal addr_of_1926_final_reg_ack_0 : boolean;
  signal type_cast_2070_inst_req_0 : boolean;
  signal addr_of_1926_final_reg_req_1 : boolean;
  signal addr_of_1926_final_reg_ack_1 : boolean;
  signal type_cast_1665_inst_ack_1 : boolean;
  signal type_cast_1665_inst_req_1 : boolean;
  signal phi_stmt_1653_req_1 : boolean;
  signal type_cast_1658_inst_ack_1 : boolean;
  signal type_cast_1658_inst_req_1 : boolean;
  signal ptr_deref_1929_store_0_req_0 : boolean;
  signal ptr_deref_1929_store_0_ack_0 : boolean;
  signal ptr_deref_1929_store_0_req_1 : boolean;
  signal ptr_deref_1929_store_0_ack_1 : boolean;
  signal type_cast_1937_inst_req_0 : boolean;
  signal type_cast_1937_inst_ack_0 : boolean;
  signal type_cast_1937_inst_req_1 : boolean;
  signal type_cast_1937_inst_ack_1 : boolean;
  signal if_stmt_1952_branch_req_0 : boolean;
  signal if_stmt_1952_branch_ack_1 : boolean;
  signal if_stmt_1952_branch_ack_0 : boolean;
  signal type_cast_1976_inst_req_0 : boolean;
  signal type_cast_1976_inst_ack_0 : boolean;
  signal type_cast_1976_inst_req_1 : boolean;
  signal type_cast_1976_inst_ack_1 : boolean;
  signal ptr_deref_1988_load_0_req_0 : boolean;
  signal ptr_deref_1988_load_0_ack_0 : boolean;
  signal ptr_deref_1988_load_0_req_1 : boolean;
  signal ptr_deref_1988_load_0_ack_1 : boolean;
  signal type_cast_2002_inst_req_0 : boolean;
  signal type_cast_2002_inst_ack_0 : boolean;
  signal type_cast_2002_inst_req_1 : boolean;
  signal type_cast_2002_inst_ack_1 : boolean;
  signal type_cast_2018_inst_req_0 : boolean;
  signal type_cast_2018_inst_ack_0 : boolean;
  signal type_cast_2018_inst_req_1 : boolean;
  signal type_cast_2018_inst_ack_1 : boolean;
  signal ptr_deref_2030_load_0_req_0 : boolean;
  signal ptr_deref_2030_load_0_ack_0 : boolean;
  signal ptr_deref_2030_load_0_req_1 : boolean;
  signal ptr_deref_2030_load_0_ack_1 : boolean;
  signal if_stmt_2048_branch_req_0 : boolean;
  signal if_stmt_2048_branch_ack_1 : boolean;
  signal if_stmt_2048_branch_ack_0 : boolean;
  signal WPIPE_Block1_complete_2078_inst_req_0 : boolean;
  signal WPIPE_Block1_complete_2078_inst_ack_0 : boolean;
  signal WPIPE_Block1_complete_2078_inst_req_1 : boolean;
  signal WPIPE_Block1_complete_2078_inst_ack_1 : boolean;
  signal phi_stmt_1659_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_B_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_B_CP_4205_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_B_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_B_CP_4205_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_B_CP_4205_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_B_CP_4205_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_B_CP_4205: Block -- control-path 
    signal zeropad3D_B_CP_4205_elements: BooleanArray(136 downto 0);
    -- 
  begin -- 
    zeropad3D_B_CP_4205_elements(0) <= zeropad3D_B_CP_4205_start;
    zeropad3D_B_CP_4205_symbol <= zeropad3D_B_CP_4205_elements(90);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1483/$entry
      -- CP-element group 0: 	 branch_block_stmt_1483/assign_stmt_1486__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1483/branch_block_stmt_1483__entry__
      -- CP-element group 0: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1483/assign_stmt_1486/$entry
      -- 
    rr_4283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(0), ack => RPIPE_Block1_starting_1485_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	136 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	97 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	100 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	104 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1483/merge_stmt_2054__exit__
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/$entry
      -- CP-element group 1: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Update/cr
      -- 
    rr_5428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(1), ack => type_cast_1665_inst_req_0); -- 
    rr_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(1), ack => type_cast_1658_inst_req_0); -- 
    cr_5479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(1), ack => type_cast_1652_inst_req_1); -- 
    rr_5474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(1), ack => type_cast_1652_inst_req_0); -- 
    cr_5433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(1), ack => type_cast_1665_inst_req_1); -- 
    cr_5456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(1), ack => type_cast_1658_inst_req_1); -- 
    zeropad3D_B_CP_4205_elements(1) <= zeropad3D_B_CP_4205_elements(136);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Sample/ra
      -- 
    ra_4284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1485_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(2)); -- 
    cr_4288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(2), ack => RPIPE_Block1_starting_1485_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: 	17 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	14 
    -- CP-element group 3: 	10 
    -- CP-element group 3: 	13 
    -- CP-element group 3: 	11 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	7 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	9 
    -- CP-element group 3:  members (129) 
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1486__exit__
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643__entry__
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1486/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1486/RPIPE_Block1_starting_1485_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_word_addrgen/root_register_ack
      -- 
    ca_4289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1485_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(3)); -- 
    cr_4383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => LOAD_pad_1511_load_0_req_1); -- 
    rr_4372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => LOAD_pad_1511_load_0_req_0); -- 
    rr_4422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1523_load_0_req_0); -- 
    cr_4433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1523_load_0_req_1); -- 
    cr_4336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1498_load_0_req_1); -- 
    cr_4355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => type_cast_1508_inst_req_1); -- 
    cr_4533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1547_load_0_req_1); -- 
    rr_4522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1547_load_0_req_0); -- 
    cr_4483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1535_load_0_req_1); -- 
    cr_4552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => type_cast_1607_inst_req_1); -- 
    rr_4472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1535_load_0_req_0); -- 
    rr_4325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(3), ack => ptr_deref_1498_load_0_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/word_access_start/word_0/ra
      -- CP-element group 4: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Sample/word_access_start/$exit
      -- 
    ra_4326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1498_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (12) 
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/word_access_complete/word_0/ca
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/ptr_deref_1498_Merge/$entry
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/ptr_deref_1498_Merge/$exit
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/ptr_deref_1498_Merge/merge_req
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/ptr_deref_1498_Merge/merge_ack
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1498_Update/$exit
      -- 
    ca_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1498_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(5)); -- 
    rr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(5), ack => type_cast_1508_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Sample/$exit
      -- 
    ra_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1508_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	3 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	18 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1508_Update/$exit
      -- 
    ca_4356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1508_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Sample/word_access_start/$exit
      -- 
    ra_4373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1511_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	3 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (12) 
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/LOAD_pad_1511_Merge/merge_ack
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/LOAD_pad_1511_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/LOAD_pad_1511_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/LOAD_pad_1511_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/LOAD_pad_1511_Update/word_access_complete/word_0/$exit
      -- 
    ca_4384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1511_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(9)); -- 
    rr_4547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(9), ack => type_cast_1607_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/word_access_start/word_0/ra
      -- CP-element group 10: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Sample/word_access_start/$exit
      -- CP-element group 10: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_sample_completed_
      -- 
    ra_4423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1523_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	18 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/word_access_complete/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/ptr_deref_1523_Merge/merge_req
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/ptr_deref_1523_Merge/merge_ack
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/word_access_complete/$exit
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/word_access_complete/word_0/ca
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/ptr_deref_1523_Merge/$entry
      -- CP-element group 11: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1523_Update/ptr_deref_1523_Merge/$exit
      -- 
    ca_4434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1523_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/word_access_start/$exit
      -- CP-element group 12: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/word_access_start/word_0/ra
      -- CP-element group 12: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Sample/$exit
      -- 
    ra_4473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1535_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	18 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/ptr_deref_1535_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/ptr_deref_1535_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/ptr_deref_1535_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1535_Update/ptr_deref_1535_Merge/merge_ack
      -- 
    ca_4484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1535_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	3 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Sample/word_access_start/word_0/ra
      -- CP-element group 14: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_sample_completed_
      -- 
    ra_4523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1547_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/ptr_deref_1547_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/ptr_deref_1547_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/ptr_deref_1547_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/ptr_deref_1547_Merge/merge_ack
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/ptr_deref_1547_update_completed_
      -- 
    ca_4534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1547_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Sample/ra
      -- 
    ra_4548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/type_cast_1607_Update/ca
      -- 
    ca_4553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(17)); -- 
    -- CP-element group 18:  join  fork  transition  place  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	11 
    -- CP-element group 18: 	7 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	91 
    -- CP-element group 18: 	92 
    -- CP-element group 18: 	93 
    -- CP-element group 18: 	95 
    -- CP-element group 18:  members (16) 
      -- CP-element group 18: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643/$exit
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/assign_stmt_1495_to_assign_stmt_1643__exit__
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1646/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1659/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/$entry
      -- CP-element group 18: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/$entry
      -- 
    cr_5399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(18), ack => type_cast_1656_inst_req_1); -- 
    rr_5394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(18), ack => type_cast_1656_inst_req_0); -- 
    zeropad3D_B_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(15) & zeropad3D_B_CP_4205_elements(17) & zeropad3D_B_CP_4205_elements(13) & zeropad3D_B_CP_4205_elements(11) & zeropad3D_B_CP_4205_elements(7);
      gj_zeropad3D_B_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	111 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Sample/ra
      -- 
    ra_4565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(19)); -- 
    -- CP-element group 20:  branch  transition  place  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	111 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (13) 
      -- CP-element group 20: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678__exit__
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679__entry__
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679_dead_link/$entry
      -- CP-element group 20: 	 branch_block_stmt_1483/R_cmp_1680_place
      -- CP-element group 20: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/$exit
      -- CP-element group 20: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679_eval_test/$entry
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679_eval_test/$exit
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679_eval_test/branch_req
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679_if_link/$entry
      -- CP-element group 20: 	 branch_block_stmt_1483/if_stmt_1679_else_link/$entry
      -- 
    ca_4570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(20)); -- 
    branch_req_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(20), ack => if_stmt_1679_branch_req_0); -- 
    -- CP-element group 21:  transition  place  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	112 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1483/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 21: 	 branch_block_stmt_1483/whilex_xbody_ifx_xthen
      -- CP-element group 21: 	 branch_block_stmt_1483/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 21: 	 branch_block_stmt_1483/if_stmt_1679_if_link/$exit
      -- CP-element group 21: 	 branch_block_stmt_1483/if_stmt_1679_if_link/if_choice_transition
      -- 
    if_choice_transition_4583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1679_branch_ack_1, ack => zeropad3D_B_CP_4205_elements(21)); -- 
    -- CP-element group 22:  merge  transition  place  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (11) 
      -- CP-element group 22: 	 branch_block_stmt_1483/merge_stmt_1685__exit__
      -- CP-element group 22: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713__entry__
      -- CP-element group 22: 	 branch_block_stmt_1483/merge_stmt_1685_PhiReqMerge
      -- CP-element group 22: 	 branch_block_stmt_1483/if_stmt_1679_else_link/$exit
      -- CP-element group 22: 	 branch_block_stmt_1483/if_stmt_1679_else_link/else_choice_transition
      -- CP-element group 22: 	 branch_block_stmt_1483/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 22: 	 branch_block_stmt_1483/merge_stmt_1685_PhiAck/dummy
      -- CP-element group 22: 	 branch_block_stmt_1483/merge_stmt_1685_PhiAck/$exit
      -- CP-element group 22: 	 branch_block_stmt_1483/merge_stmt_1685_PhiAck/$entry
      -- CP-element group 22: 	 branch_block_stmt_1483/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 22: 	 branch_block_stmt_1483/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- 
    else_choice_transition_4587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1679_branch_ack_0, ack => zeropad3D_B_CP_4205_elements(22)); -- 
    -- CP-element group 23:  join  fork  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (27) 
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_address_calculated
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_word_address_calculated
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_root_address_calculated
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_address_resized
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_addr_resize/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_addr_resize/$exit
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_addr_resize/base_resize_req
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_addr_resize/base_resize_ack
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_plus_offset/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_plus_offset/$exit
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_plus_offset/sum_rename_req
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_base_plus_offset/sum_rename_ack
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_word_addrgen/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_word_addrgen/$exit
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_word_addrgen/root_register_req
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_word_addrgen/root_register_ack
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/word_access_start/word_0/rr
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/word_access_complete/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/word_access_complete/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/word_access_complete/word_0/cr
      -- 
    cr_4636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(23), ack => ptr_deref_1696_load_0_req_1); -- 
    rr_4625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(23), ack => ptr_deref_1696_load_0_req_0); -- 
    zeropad3D_B_CP_4205_elements(23) <= zeropad3D_B_CP_4205_elements(22);
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Sample/word_access_start/word_0/ra
      -- 
    ra_4626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1696_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(24)); -- 
    -- CP-element group 25:  branch  transition  place  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (19) 
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713__exit__
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714__entry__
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/$exit
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/ptr_deref_1696_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/ptr_deref_1696_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/ptr_deref_1696_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_1483/assign_stmt_1693_to_assign_stmt_1713/ptr_deref_1696_Update/ptr_deref_1696_Merge/merge_ack
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714_dead_link/$entry
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714_eval_test/$entry
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714_eval_test/$exit
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714_eval_test/branch_req
      -- CP-element group 25: 	 branch_block_stmt_1483/R_cmp50_1715_place
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714_if_link/$entry
      -- CP-element group 25: 	 branch_block_stmt_1483/if_stmt_1714_else_link/$entry
      -- 
    ca_4637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1696_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(25)); -- 
    branch_req_4650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(25), ack => if_stmt_1714_branch_req_0); -- 
    -- CP-element group 26:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (18) 
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732__entry__
      -- CP-element group 26: 	 branch_block_stmt_1483/merge_stmt_1720__exit__
      -- CP-element group 26: 	 branch_block_stmt_1483/merge_stmt_1720_PhiReqMerge
      -- CP-element group 26: 	 branch_block_stmt_1483/if_stmt_1714_if_link/$exit
      -- CP-element group 26: 	 branch_block_stmt_1483/if_stmt_1714_if_link/if_choice_transition
      -- CP-element group 26: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse52
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/$entry
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_1483/merge_stmt_1720_PhiAck/dummy
      -- CP-element group 26: 	 branch_block_stmt_1483/merge_stmt_1720_PhiAck/$exit
      -- CP-element group 26: 	 branch_block_stmt_1483/merge_stmt_1720_PhiAck/$entry
      -- CP-element group 26: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse52_PhiReq/$exit
      -- CP-element group 26: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse52_PhiReq/$entry
      -- 
    if_choice_transition_4655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1714_branch_ack_1, ack => zeropad3D_B_CP_4205_elements(26)); -- 
    rr_4672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(26), ack => type_cast_1724_inst_req_0); -- 
    cr_4677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(26), ack => type_cast_1724_inst_req_1); -- 
    -- CP-element group 27:  transition  place  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	112 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- CP-element group 27: 	 branch_block_stmt_1483/if_stmt_1714_else_link/$exit
      -- CP-element group 27: 	 branch_block_stmt_1483/if_stmt_1714_else_link/else_choice_transition
      -- CP-element group 27: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse_ifx_xthen
      -- 
    else_choice_transition_4659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1714_branch_ack_0, ack => zeropad3D_B_CP_4205_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Sample/ra
      -- 
    ra_4673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(28)); -- 
    -- CP-element group 29:  branch  transition  place  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (13) 
      -- CP-element group 29: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732__exit__
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733__entry__
      -- CP-element group 29: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/$exit
      -- CP-element group 29: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1483/assign_stmt_1725_to_assign_stmt_1732/type_cast_1724_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733_dead_link/$entry
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733_eval_test/$entry
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733_eval_test/$exit
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733_eval_test/branch_req
      -- CP-element group 29: 	 branch_block_stmt_1483/R_cmp57_1734_place
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733_if_link/$entry
      -- CP-element group 29: 	 branch_block_stmt_1483/if_stmt_1733_else_link/$entry
      -- 
    ca_4678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(29)); -- 
    branch_req_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(29), ack => if_stmt_1733_branch_req_0); -- 
    -- CP-element group 30:  transition  place  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	112 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse52_ifx_xthen_PhiReq/$exit
      -- CP-element group 30: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse52_ifx_xthen_PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_1483/if_stmt_1733_if_link/$exit
      -- CP-element group 30: 	 branch_block_stmt_1483/if_stmt_1733_if_link/if_choice_transition
      -- CP-element group 30: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse52_ifx_xthen
      -- 
    if_choice_transition_4691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1733_branch_ack_1, ack => zeropad3D_B_CP_4205_elements(30)); -- 
    -- CP-element group 31:  merge  transition  place  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (11) 
      -- CP-element group 31: 	 branch_block_stmt_1483/merge_stmt_1739__exit__
      -- CP-element group 31: 	 branch_block_stmt_1483/merge_stmt_1739_PhiReqMerge
      -- CP-element group 31: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761__entry__
      -- CP-element group 31: 	 branch_block_stmt_1483/if_stmt_1733_else_link/$exit
      -- CP-element group 31: 	 branch_block_stmt_1483/if_stmt_1733_else_link/else_choice_transition
      -- CP-element group 31: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse52_lorx_xlhsx_xfalse59
      -- CP-element group 31: 	 branch_block_stmt_1483/merge_stmt_1739_PhiAck/dummy
      -- CP-element group 31: 	 branch_block_stmt_1483/merge_stmt_1739_PhiAck/$exit
      -- CP-element group 31: 	 branch_block_stmt_1483/merge_stmt_1739_PhiAck/$entry
      -- CP-element group 31: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse52_lorx_xlhsx_xfalse59_PhiReq/$exit
      -- CP-element group 31: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse52_lorx_xlhsx_xfalse59_PhiReq/$entry
      -- 
    else_choice_transition_4695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1733_branch_ack_0, ack => zeropad3D_B_CP_4205_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (27) 
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_address_calculated
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_word_address_calculated
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_root_address_calculated
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_address_resized
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_addr_resize/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_addr_resize/$exit
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_addr_resize/base_resize_req
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_addr_resize/base_resize_ack
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_plus_offset/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_plus_offset/$exit
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_plus_offset/sum_rename_req
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_base_plus_offset/sum_rename_ack
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_word_addrgen/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_word_addrgen/$exit
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_word_addrgen/root_register_req
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_word_addrgen/root_register_ack
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/word_access_start/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/word_access_start/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/word_access_start/word_0/rr
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/word_access_complete/word_0/cr
      -- 
    cr_4744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(32), ack => ptr_deref_1750_load_0_req_1); -- 
    rr_4733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(32), ack => ptr_deref_1750_load_0_req_0); -- 
    zeropad3D_B_CP_4205_elements(32) <= zeropad3D_B_CP_4205_elements(31);
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Sample/word_access_start/word_0/ra
      -- 
    ra_4734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1750_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (19) 
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761__exit__
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762__entry__
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/$exit
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/word_access_complete/word_0/ca
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/ptr_deref_1750_Merge/$entry
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/ptr_deref_1750_Merge/$exit
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/ptr_deref_1750_Merge/merge_req
      -- CP-element group 34: 	 branch_block_stmt_1483/assign_stmt_1747_to_assign_stmt_1761/ptr_deref_1750_Update/ptr_deref_1750_Merge/merge_ack
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762_eval_test/branch_req
      -- CP-element group 34: 	 branch_block_stmt_1483/R_cmp66_1763_place
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1483/if_stmt_1762_else_link/$entry
      -- 
    ca_4745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1750_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(34)); -- 
    branch_req_4758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(34), ack => if_stmt_1762_branch_req_0); -- 
    -- CP-element group 35:  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	51 
    -- CP-element group 35: 	52 
    -- CP-element group 35: 	54 
    -- CP-element group 35: 	56 
    -- CP-element group 35: 	58 
    -- CP-element group 35: 	60 
    -- CP-element group 35: 	62 
    -- CP-element group 35: 	64 
    -- CP-element group 35: 	66 
    -- CP-element group 35: 	69 
    -- CP-element group 35:  members (46) 
      -- CP-element group 35: 	 branch_block_stmt_1483/merge_stmt_1826__exit__
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931__entry__
      -- CP-element group 35: 	 branch_block_stmt_1483/merge_stmt_1826_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_1483/if_stmt_1762_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_1483/if_stmt_1762_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse59_ifx_xelse
      -- CP-element group 35: 	 branch_block_stmt_1483/merge_stmt_1826_PhiAck/dummy
      -- CP-element group 35: 	 branch_block_stmt_1483/merge_stmt_1826_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/merge_stmt_1826_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse59_ifx_xelse_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_update_start
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Update/req
      -- CP-element group 35: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse59_ifx_xelse_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_complete/req
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/word_access_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/word_access_complete/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/word_access_complete/word_0/cr
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_update_start
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Update/req
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_complete/req
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/word_access_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/word_access_complete/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/word_access_complete/word_0/cr
      -- 
    if_choice_transition_4763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1762_branch_ack_1, ack => zeropad3D_B_CP_4205_elements(35)); -- 
    rr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => type_cast_1830_inst_req_0); -- 
    cr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => type_cast_1830_inst_req_1); -- 
    cr_4940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => type_cast_1894_inst_req_1); -- 
    req_4971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => array_obj_ref_1900_index_offset_req_1); -- 
    req_4986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => addr_of_1901_final_reg_req_1); -- 
    cr_5031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => ptr_deref_1905_load_0_req_1); -- 
    cr_5050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => type_cast_1919_inst_req_1); -- 
    req_5081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => array_obj_ref_1925_index_offset_req_1); -- 
    req_5096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => addr_of_1926_final_reg_req_1); -- 
    cr_5146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(35), ack => ptr_deref_1929_store_0_req_1); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	112 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse59_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse59_ifx_xthen_PhiReq/$exit
      -- CP-element group 36: 	 branch_block_stmt_1483/if_stmt_1762_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_1483/if_stmt_1762_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_1483/lorx_xlhsx_xfalse59_ifx_xthen
      -- 
    else_choice_transition_4767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1762_branch_ack_0, ack => zeropad3D_B_CP_4205_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	112 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Sample/ra
      -- 
    ra_4781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	112 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Update/ca
      -- 
    ca_4786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	112 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Sample/ra
      -- 
    ra_4795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1777_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	112 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Update/ca
      -- 
    ca_4800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1777_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Sample/rr
      -- 
    rr_4808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(41), ack => type_cast_1811_inst_req_0); -- 
    zeropad3D_B_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(40) & zeropad3D_B_CP_4205_elements(38);
      gj_zeropad3D_B_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Sample/ra
      -- 
    ra_4809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1811_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	112 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (16) 
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Sample/req
      -- 
    ca_4814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1811_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(43)); -- 
    req_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(43), ack => array_obj_ref_1817_index_offset_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Sample/ack
      -- 
    ack_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1817_index_offset_ack_0, ack => zeropad3D_B_CP_4205_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	112 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (11) 
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_offset_calculated
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_request/$entry
      -- CP-element group 45: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_request/req
      -- 
    ack_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1817_index_offset_ack_1, ack => zeropad3D_B_CP_4205_elements(45)); -- 
    req_4854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(45), ack => addr_of_1818_final_reg_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_request/$exit
      -- CP-element group 46: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_request/ack
      -- 
    ack_4855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1818_final_reg_ack_0, ack => zeropad3D_B_CP_4205_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	112 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (28) 
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_complete/ack
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_word_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_address_resized
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_addr_resize/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_addr_resize/$exit
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_addr_resize/base_resize_req
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_addr_resize/base_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_word_addrgen/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_word_addrgen/$exit
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_word_addrgen/root_register_req
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_word_addrgen/root_register_ack
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/ptr_deref_1821_Split/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/ptr_deref_1821_Split/$exit
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/ptr_deref_1821_Split/split_req
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/ptr_deref_1821_Split/split_ack
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/word_access_start/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/word_access_start/word_0/$entry
      -- CP-element group 47: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/word_access_start/word_0/rr
      -- 
    ack_4860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1818_final_reg_ack_1, ack => zeropad3D_B_CP_4205_elements(47)); -- 
    rr_4898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(47), ack => ptr_deref_1821_store_0_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/word_access_start/$exit
      -- CP-element group 48: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Sample/word_access_start/word_0/ra
      -- 
    ra_4899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1821_store_0_ack_0, ack => zeropad3D_B_CP_4205_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	112 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/word_access_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/word_access_complete/word_0/ca
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1821_store_0_ack_1, ack => zeropad3D_B_CP_4205_elements(49)); -- 
    -- CP-element group 50:  join  transition  place  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	44 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	113 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824__exit__
      -- CP-element group 50: 	 branch_block_stmt_1483/ifx_xthen_ifx_xend
      -- CP-element group 50: 	 branch_block_stmt_1483/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 50: 	 branch_block_stmt_1483/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/$exit
      -- 
    zeropad3D_B_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(49) & zeropad3D_B_CP_4205_elements(44);
      gj_zeropad3D_B_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	35 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Sample/ra
      -- 
    ra_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	35 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	61 
    -- CP-element group 52:  members (9) 
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1830_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Sample/rr
      -- 
    ca_4927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(52)); -- 
    rr_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(52), ack => type_cast_1894_inst_req_0); -- 
    rr_5045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(52), ack => type_cast_1919_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Sample/ra
      -- 
    ra_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	35 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (16) 
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1894_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_resized_1
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_scaled_1
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_computed_1
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_resize_1/$entry
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_resize_1/$exit
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_resize_1/index_resize_req
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_resize_1/index_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_scale_1/$entry
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_scale_1/$exit
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_scale_1/scale_rename_req
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_index_scale_1/scale_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Sample/req
      -- 
    ca_4941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(54)); -- 
    req_4966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(54), ack => array_obj_ref_1900_index_offset_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	70 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_sample_complete
      -- CP-element group 55: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Sample/ack
      -- 
    ack_4967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1900_index_offset_ack_0, ack => zeropad3D_B_CP_4205_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	35 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (11) 
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_offset_calculated
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_final_index_sum_regn_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1900_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_request/$entry
      -- CP-element group 56: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_request/req
      -- 
    ack_4972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1900_index_offset_ack_1, ack => zeropad3D_B_CP_4205_elements(56)); -- 
    req_4981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(56), ack => addr_of_1901_final_reg_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_request/$exit
      -- CP-element group 57: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_request/ack
      -- 
    ack_4982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1901_final_reg_ack_0, ack => zeropad3D_B_CP_4205_elements(57)); -- 
    -- CP-element group 58:  join  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	35 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1901_complete/ack
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/word_access_start/word_0/rr
      -- 
    ack_4987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1901_final_reg_ack_1, ack => zeropad3D_B_CP_4205_elements(58)); -- 
    rr_5020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(58), ack => ptr_deref_1905_load_0_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Sample/word_access_start/word_0/ra
      -- 
    ra_5021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	35 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	67 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/ptr_deref_1905_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/ptr_deref_1905_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_ack
      -- 
    ca_5032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	52 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Sample/ra
      -- 
    ra_5046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	35 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (16) 
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/type_cast_1919_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_resized_1
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_scaled_1
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_computed_1
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_resize_1/$entry
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_resize_1/$exit
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_resize_1/index_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_resize_1/index_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_scale_1/$entry
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_scale_1/$exit
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_scale_1/scale_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_index_scale_1/scale_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Sample/req
      -- 
    ca_5051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(62)); -- 
    req_5076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(62), ack => array_obj_ref_1925_index_offset_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	70 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_sample_complete
      -- CP-element group 63: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Sample/ack
      -- 
    ack_5077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1925_index_offset_ack_0, ack => zeropad3D_B_CP_4205_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	35 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (11) 
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_offset_calculated
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_final_index_sum_regn_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/array_obj_ref_1925_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_request/$entry
      -- CP-element group 64: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_request/req
      -- 
    ack_5082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1925_index_offset_ack_1, ack => zeropad3D_B_CP_4205_elements(64)); -- 
    req_5091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(64), ack => addr_of_1926_final_reg_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_request/$exit
      -- CP-element group 65: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_request/ack
      -- 
    ack_5092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1926_final_reg_ack_0, ack => zeropad3D_B_CP_4205_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	35 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (19) 
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/addr_of_1926_complete/ack
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_word_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_root_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_address_resized
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_addr_resize/$entry
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_addr_resize/$exit
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_addr_resize/base_resize_req
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_addr_resize/base_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_plus_offset/$entry
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_plus_offset/$exit
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_plus_offset/sum_rename_req
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_base_plus_offset/sum_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_word_addrgen/$entry
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_word_addrgen/$exit
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_word_addrgen/root_register_req
      -- CP-element group 66: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_word_addrgen/root_register_ack
      -- 
    ack_5097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1926_final_reg_ack_1, ack => zeropad3D_B_CP_4205_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	60 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/ptr_deref_1929_Split/$entry
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/ptr_deref_1929_Split/$exit
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/ptr_deref_1929_Split/split_req
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/ptr_deref_1929_Split/split_ack
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/word_access_start/$entry
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/word_access_start/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/word_access_start/word_0/rr
      -- 
    rr_5135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(67), ack => ptr_deref_1929_store_0_req_0); -- 
    zeropad3D_B_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(60) & zeropad3D_B_CP_4205_elements(66);
      gj_zeropad3D_B_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/word_access_start/$exit
      -- CP-element group 68: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/word_access_start/word_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Sample/word_access_start/word_0/ra
      -- 
    ra_5136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1929_store_0_ack_0, ack => zeropad3D_B_CP_4205_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	35 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/word_access_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/word_access_complete/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/ptr_deref_1929_Update/word_access_complete/word_0/ca
      -- 
    ca_5147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1929_store_0_ack_1, ack => zeropad3D_B_CP_4205_elements(69)); -- 
    -- CP-element group 70:  join  transition  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	55 
    -- CP-element group 70: 	63 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	113 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1483/ifx_xelse_ifx_xend
      -- CP-element group 70: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931__exit__
      -- CP-element group 70: 	 branch_block_stmt_1483/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1483/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1483/assign_stmt_1831_to_assign_stmt_1931/$exit
      -- 
    zeropad3D_B_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(55) & zeropad3D_B_CP_4205_elements(63) & zeropad3D_B_CP_4205_elements(69);
      gj_zeropad3D_B_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	113 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Sample/ra
      -- 
    ra_5159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(71)); -- 
    -- CP-element group 72:  branch  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	113 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (13) 
      -- CP-element group 72: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951__exit__
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952__entry__
      -- CP-element group 72: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/$exit
      -- CP-element group 72: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952_dead_link/$entry
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952_eval_test/$entry
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952_eval_test/$exit
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952_eval_test/branch_req
      -- CP-element group 72: 	 branch_block_stmt_1483/R_cmp135_1953_place
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952_if_link/$entry
      -- CP-element group 72: 	 branch_block_stmt_1483/if_stmt_1952_else_link/$entry
      -- 
    ca_5164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(72)); -- 
    branch_req_5172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(72), ack => if_stmt_1952_branch_req_0); -- 
    -- CP-element group 73:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	122 
    -- CP-element group 73: 	123 
    -- CP-element group 73: 	125 
    -- CP-element group 73: 	126 
    -- CP-element group 73: 	128 
    -- CP-element group 73: 	129 
    -- CP-element group 73:  members (40) 
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xend_ifx_xthen137_PhiReq/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/merge_stmt_1958__exit__
      -- CP-element group 73: 	 branch_block_stmt_1483/assign_stmt_1964__entry__
      -- CP-element group 73: 	 branch_block_stmt_1483/assign_stmt_1964__exit__
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Update/cr
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/cr
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Update/cr
      -- CP-element group 73: 	 branch_block_stmt_1483/merge_stmt_1958_PhiAck/dummy
      -- CP-element group 73: 	 branch_block_stmt_1483/merge_stmt_1958_PhiAck/$exit
      -- CP-element group 73: 	 branch_block_stmt_1483/merge_stmt_1958_PhiAck/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_1483/merge_stmt_1958_PhiReqMerge
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xend_ifx_xthen137_PhiReq/$exit
      -- CP-element group 73: 	 branch_block_stmt_1483/if_stmt_1952_if_link/$exit
      -- CP-element group 73: 	 branch_block_stmt_1483/if_stmt_1952_if_link/if_choice_transition
      -- CP-element group 73: 	 branch_block_stmt_1483/ifx_xend_ifx_xthen137
      -- CP-element group 73: 	 branch_block_stmt_1483/assign_stmt_1964/$entry
      -- CP-element group 73: 	 branch_block_stmt_1483/assign_stmt_1964/$exit
      -- 
    if_choice_transition_5177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1952_branch_ack_1, ack => zeropad3D_B_CP_4205_elements(73)); -- 
    cr_5715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(73), ack => type_cast_2060_inst_req_1); -- 
    cr_5669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(73), ack => type_cast_2064_inst_req_1); -- 
    rr_5664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(73), ack => type_cast_2064_inst_req_0); -- 
    rr_5710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(73), ack => type_cast_2060_inst_req_0); -- 
    cr_5692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(73), ack => type_cast_2070_inst_req_1); -- 
    rr_5687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(73), ack => type_cast_2070_inst_req_0); -- 
    -- CP-element group 74:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74: 	77 
    -- CP-element group 74: 	78 
    -- CP-element group 74: 	81 
    -- CP-element group 74: 	83 
    -- CP-element group 74: 	84 
    -- CP-element group 74: 	85 
    -- CP-element group 74:  members (76) 
      -- CP-element group 74: 	 branch_block_stmt_1483/merge_stmt_1966__exit__
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047__entry__
      -- CP-element group 74: 	 branch_block_stmt_1483/merge_stmt_1966_PhiAck/dummy
      -- CP-element group 74: 	 branch_block_stmt_1483/merge_stmt_1966_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/merge_stmt_1966_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/merge_stmt_1966_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_1483/ifx_xend_ifx_xelse142_PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/ifx_xend_ifx_xelse142_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/if_stmt_1952_else_link/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/if_stmt_1952_else_link/else_choice_transition
      -- CP-element group 74: 	 branch_block_stmt_1483/ifx_xend_ifx_xelse142
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_address_calculated
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_word_address_calculated
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_root_address_calculated
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_address_resized
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_addr_resize/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_addr_resize/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_addr_resize/base_resize_req
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_addr_resize/base_resize_ack
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_plus_offset/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_plus_offset/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_plus_offset/sum_rename_req
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_base_plus_offset/sum_rename_ack
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_word_addrgen/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_word_addrgen/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_word_addrgen/root_register_req
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_word_addrgen/root_register_ack
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/word_access_complete/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/word_access_complete/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/word_access_complete/word_0/cr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_address_calculated
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_word_address_calculated
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_root_address_calculated
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_address_resized
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_addr_resize/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_addr_resize/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_addr_resize/base_resize_req
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_addr_resize/base_resize_ack
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_plus_offset/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_plus_offset/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_plus_offset/sum_rename_req
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_base_plus_offset/sum_rename_ack
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_word_addrgen/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_word_addrgen/$exit
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_word_addrgen/root_register_req
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_word_addrgen/root_register_ack
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/word_access_complete/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/word_access_complete/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1952_branch_ack_0, ack => zeropad3D_B_CP_4205_elements(74)); -- 
    rr_5197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => type_cast_1976_inst_req_0); -- 
    cr_5202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => type_cast_1976_inst_req_1); -- 
    rr_5236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => ptr_deref_1988_load_0_req_0); -- 
    cr_5247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => ptr_deref_1988_load_0_req_1); -- 
    cr_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => type_cast_2002_inst_req_1); -- 
    cr_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => type_cast_2018_inst_req_1); -- 
    rr_5314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => ptr_deref_2030_load_0_req_0); -- 
    cr_5325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(74), ack => ptr_deref_2030_load_0_req_1); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Sample/ra
      -- 
    ra_5198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	79 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_1976_Update/ca
      -- 
    ca_5203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/word_access_start/$exit
      -- CP-element group 77: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/word_access_start/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Sample/word_access_start/word_0/ra
      -- 
    ra_5237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/word_access_complete/$exit
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/word_access_complete/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/word_access_complete/word_0/ca
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/ptr_deref_1988_Merge/$entry
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/ptr_deref_1988_Merge/$exit
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/ptr_deref_1988_Merge/merge_req
      -- CP-element group 78: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_1988_Update/ptr_deref_1988_Merge/merge_ack
      -- 
    ca_5248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	76 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Sample/rr
      -- 
    rr_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(79), ack => type_cast_2002_inst_req_0); -- 
    zeropad3D_B_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(76) & zeropad3D_B_CP_4205_elements(78);
      gj_zeropad3D_B_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Sample/ra
      -- 
    ra_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	74 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2002_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Sample/rr
      -- 
    ca_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(81)); -- 
    rr_5275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(81), ack => type_cast_2018_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Sample/ra
      -- 
    ra_5276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	74 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/type_cast_2018_Update/ca
      -- 
    ca_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	74 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/word_access_start/$exit
      -- CP-element group 84: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Sample/word_access_start/word_0/ra
      -- 
    ra_5315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2030_load_0_ack_0, ack => zeropad3D_B_CP_4205_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	74 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/word_access_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/word_access_complete/word_0/ca
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/ptr_deref_2030_Merge/$entry
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/ptr_deref_2030_Merge/$exit
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/ptr_deref_2030_Merge/merge_req
      -- CP-element group 85: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/ptr_deref_2030_Update/ptr_deref_2030_Merge/merge_ack
      -- 
    ca_5326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2030_load_0_ack_1, ack => zeropad3D_B_CP_4205_elements(85)); -- 
    -- CP-element group 86:  branch  join  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (10) 
      -- CP-element group 86: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047__exit__
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048__entry__
      -- CP-element group 86: 	 branch_block_stmt_1483/assign_stmt_1972_to_assign_stmt_2047/$exit
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_1483/R_cmp165_2049_place
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_1483/if_stmt_2048_else_link/$entry
      -- 
    branch_req_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(86), ack => if_stmt_2048_branch_req_0); -- 
    zeropad3D_B_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(83) & zeropad3D_B_CP_4205_elements(85);
      gj_zeropad3D_B_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (15) 
      -- CP-element group 87: 	 branch_block_stmt_1483/ifx_xelse142_whilex_xend_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_1483/assign_stmt_2080__entry__
      -- CP-element group 87: 	 branch_block_stmt_1483/merge_stmt_2076__exit__
      -- CP-element group 87: 	 branch_block_stmt_1483/merge_stmt_2076_PhiAck/dummy
      -- CP-element group 87: 	 branch_block_stmt_1483/merge_stmt_2076_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_1483/merge_stmt_2076_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_1483/merge_stmt_2076_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1483/ifx_xelse142_whilex_xend_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_1483/if_stmt_2048_if_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_1483/if_stmt_2048_if_link/if_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_1483/ifx_xelse142_whilex_xend
      -- CP-element group 87: 	 branch_block_stmt_1483/assign_stmt_2080/$entry
      -- CP-element group 87: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Sample/req
      -- 
    if_choice_transition_5344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2048_branch_ack_1, ack => zeropad3D_B_CP_4205_elements(87)); -- 
    req_5361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(87), ack => WPIPE_Block1_complete_2078_inst_req_0); -- 
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	114 
    -- CP-element group 88: 	115 
    -- CP-element group 88: 	117 
    -- CP-element group 88: 	118 
    -- CP-element group 88: 	119 
    -- CP-element group 88:  members (22) 
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2067/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/$entry
      -- CP-element group 88: 	 branch_block_stmt_1483/if_stmt_2048_else_link/$exit
      -- CP-element group 88: 	 branch_block_stmt_1483/if_stmt_2048_else_link/else_choice_transition
      -- CP-element group 88: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173
      -- 
    else_choice_transition_5348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2048_branch_ack_0, ack => zeropad3D_B_CP_4205_elements(88)); -- 
    cr_5612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(88), ack => type_cast_2066_inst_req_1); -- 
    rr_5607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(88), ack => type_cast_2066_inst_req_0); -- 
    cr_5643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(88), ack => type_cast_2058_inst_req_1); -- 
    rr_5638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(88), ack => type_cast_2058_inst_req_0); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Update/req
      -- 
    ack_5362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_complete_2078_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(89)); -- 
    req_5366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(89), ack => WPIPE_Block1_complete_2078_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (16) 
      -- CP-element group 90: 	 $exit
      -- CP-element group 90: 	 branch_block_stmt_1483/branch_block_stmt_1483__exit__
      -- CP-element group 90: 	 branch_block_stmt_1483/$exit
      -- CP-element group 90: 	 branch_block_stmt_1483/merge_stmt_2082__exit__
      -- CP-element group 90: 	 branch_block_stmt_1483/return__
      -- CP-element group 90: 	 branch_block_stmt_1483/assign_stmt_2080__exit__
      -- CP-element group 90: 	 branch_block_stmt_1483/merge_stmt_2082_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_1483/return___PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_1483/return___PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_1483/merge_stmt_2082_PhiAck/dummy
      -- CP-element group 90: 	 branch_block_stmt_1483/merge_stmt_2082_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_1483/merge_stmt_2082_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_1483/assign_stmt_2080/$exit
      -- CP-element group 90: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1483/assign_stmt_2080/WPIPE_Block1_complete_2078_Update/ack
      -- 
    ack_5367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_complete_2078_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(90)); -- 
    -- CP-element group 91:  transition  output  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	18 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	96 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1659/$exit
      -- CP-element group 91: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1663_konst_delay_trans
      -- CP-element group 91: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_req
      -- 
    phi_stmt_1659_req_5378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1659_req_5378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(91), ack => phi_stmt_1659_req_0); -- 
    -- Element group zeropad3D_B_CP_4205_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_4205_elements(18), ack => zeropad3D_B_CP_4205_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Sample/$exit
      -- 
    ra_5395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1656_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	18 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Update/ca
      -- CP-element group 93: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/Update/$exit
      -- 
    ca_5400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1656_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_req
      -- CP-element group 94: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/$exit
      -- CP-element group 94: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/$exit
      -- CP-element group 94: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1656/SplitProtocol/$exit
      -- 
    phi_stmt_1653_req_5401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1653_req_5401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(94), ack => phi_stmt_1653_req_0); -- 
    zeropad3D_B_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(92) & zeropad3D_B_CP_4205_elements(93);
      gj_zeropad3D_B_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  output  delay-element  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	18 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_req
      -- CP-element group 95: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1650_konst_delay_trans
      -- CP-element group 95: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/phi_stmt_1646/$exit
      -- 
    phi_stmt_1646_req_5409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1646_req_5409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(95), ack => phi_stmt_1646_req_0); -- 
    -- Element group zeropad3D_B_CP_4205_elements(95) is a control-delay.
    cp_element_95_delay: control_delay_element  generic map(name => " 95_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_4205_elements(18), ack => zeropad3D_B_CP_4205_elements(95), clk => clk, reset =>reset);
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	91 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	107 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1483/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(91) & zeropad3D_B_CP_4205_elements(94) & zeropad3D_B_CP_4205_elements(95);
      gj_zeropad3D_B_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	1 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Sample/$exit
      -- 
    ra_5429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Update/ca
      -- CP-element group 98: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/Update/$exit
      -- 
    ca_5434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	106 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/SplitProtocol/$exit
      -- CP-element group 99: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/type_cast_1665/$exit
      -- CP-element group 99: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/$exit
      -- CP-element group 99: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1659/phi_stmt_1659_req
      -- 
    phi_stmt_1659_req_5435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1659_req_5435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(99), ack => phi_stmt_1659_req_1); -- 
    zeropad3D_B_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(97) & zeropad3D_B_CP_4205_elements(98);
      gj_zeropad3D_B_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Sample/$exit
      -- 
    ra_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/Update/ca
      -- 
    ca_5457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(101)); -- 
    -- CP-element group 102:  join  transition  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	106 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/$exit
      -- CP-element group 102: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/SplitProtocol/$exit
      -- CP-element group 102: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_sources/type_cast_1658/$exit
      -- CP-element group 102: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/$exit
      -- CP-element group 102: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1653/phi_stmt_1653_req
      -- 
    phi_stmt_1653_req_5458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1653_req_5458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(102), ack => phi_stmt_1653_req_1); -- 
    zeropad3D_B_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(100) & zeropad3D_B_CP_4205_elements(101);
      gj_zeropad3D_B_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Sample/$exit
      -- 
    ra_5475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1652_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	1 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/Update/$exit
      -- 
    ca_5480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1652_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_req
      -- CP-element group 105: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/type_cast_1652/$exit
      -- CP-element group 105: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/phi_stmt_1646_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/phi_stmt_1646/$exit
      -- 
    phi_stmt_1646_req_5481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1646_req_5481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(105), ack => phi_stmt_1646_req_1); -- 
    zeropad3D_B_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(103) & zeropad3D_B_CP_4205_elements(104);
      gj_zeropad3D_B_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	99 
    -- CP-element group 106: 	102 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1483/ifx_xend173_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(99) & zeropad3D_B_CP_4205_elements(102) & zeropad3D_B_CP_4205_elements(105);
      gj_zeropad3D_B_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  merge  fork  transition  place  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	96 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	109 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1483/merge_stmt_1645_PhiReqMerge
      -- CP-element group 107: 	 branch_block_stmt_1483/merge_stmt_1645_PhiAck/$entry
      -- 
    zeropad3D_B_CP_4205_elements(107) <= OrReduce(zeropad3D_B_CP_4205_elements(96) & zeropad3D_B_CP_4205_elements(106));
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1483/merge_stmt_1645_PhiAck/phi_stmt_1646_ack
      -- 
    phi_stmt_1646_ack_5486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1646_ack_0, ack => zeropad3D_B_CP_4205_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1483/merge_stmt_1645_PhiAck/phi_stmt_1653_ack
      -- 
    phi_stmt_1653_ack_5487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1653_ack_0, ack => zeropad3D_B_CP_4205_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1483/merge_stmt_1645_PhiAck/phi_stmt_1659_ack
      -- 
    phi_stmt_1659_ack_5488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1659_ack_0, ack => zeropad3D_B_CP_4205_elements(110)); -- 
    -- CP-element group 111:  join  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	19 
    -- CP-element group 111: 	20 
    -- CP-element group 111:  members (10) 
      -- CP-element group 111: 	 branch_block_stmt_1483/merge_stmt_1645__exit__
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678__entry__
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/$entry
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1483/assign_stmt_1671_to_assign_stmt_1678/type_cast_1670_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_1483/merge_stmt_1645_PhiAck/$exit
      -- 
    rr_4564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(111), ack => type_cast_1670_inst_req_0); -- 
    cr_4569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(111), ack => type_cast_1670_inst_req_1); -- 
    zeropad3D_B_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(108) & zeropad3D_B_CP_4205_elements(109) & zeropad3D_B_CP_4205_elements(110);
      gj_zeropad3D_B_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  merge  fork  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	27 
    -- CP-element group 112: 	21 
    -- CP-element group 112: 	30 
    -- CP-element group 112: 	36 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	49 
    -- CP-element group 112: 	47 
    -- CP-element group 112: 	45 
    -- CP-element group 112: 	39 
    -- CP-element group 112: 	40 
    -- CP-element group 112: 	43 
    -- CP-element group 112: 	37 
    -- CP-element group 112: 	38 
    -- CP-element group 112:  members (33) 
      -- CP-element group 112: 	 branch_block_stmt_1483/merge_stmt_1768__exit__
      -- CP-element group 112: 	 branch_block_stmt_1483/merge_stmt_1768_PhiAck/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824__entry__
      -- CP-element group 112: 	 branch_block_stmt_1483/merge_stmt_1768_PhiAck/$exit
      -- CP-element group 112: 	 branch_block_stmt_1483/merge_stmt_1768_PhiReqMerge
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1772_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1777_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/type_cast_1811_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_update_start
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/array_obj_ref_1817_final_index_sum_regn_Update/req
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_complete/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/addr_of_1818_complete/req
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/word_access_complete/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/word_access_complete/word_0/$entry
      -- CP-element group 112: 	 branch_block_stmt_1483/assign_stmt_1773_to_assign_stmt_1824/ptr_deref_1821_Update/word_access_complete/word_0/cr
      -- CP-element group 112: 	 branch_block_stmt_1483/merge_stmt_1768_PhiAck/dummy
      -- 
    rr_4780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => type_cast_1772_inst_req_0); -- 
    cr_4785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => type_cast_1772_inst_req_1); -- 
    rr_4794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => type_cast_1777_inst_req_0); -- 
    cr_4799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => type_cast_1777_inst_req_1); -- 
    cr_4813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => type_cast_1811_inst_req_1); -- 
    req_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => array_obj_ref_1817_index_offset_req_1); -- 
    req_4859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => addr_of_1818_final_reg_req_1); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(112), ack => ptr_deref_1821_store_0_req_1); -- 
    zeropad3D_B_CP_4205_elements(112) <= OrReduce(zeropad3D_B_CP_4205_elements(27) & zeropad3D_B_CP_4205_elements(21) & zeropad3D_B_CP_4205_elements(30) & zeropad3D_B_CP_4205_elements(36));
    -- CP-element group 113:  merge  fork  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	50 
    -- CP-element group 113: 	70 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	71 
    -- CP-element group 113: 	72 
    -- CP-element group 113:  members (13) 
      -- CP-element group 113: 	 branch_block_stmt_1483/merge_stmt_1933__exit__
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951__entry__
      -- CP-element group 113: 	 branch_block_stmt_1483/merge_stmt_1933_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_1483/merge_stmt_1933_PhiAck/$exit
      -- CP-element group 113: 	 branch_block_stmt_1483/merge_stmt_1933_PhiAck/$entry
      -- CP-element group 113: 	 branch_block_stmt_1483/merge_stmt_1933_PhiAck/dummy
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/$entry
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1483/assign_stmt_1938_to_assign_stmt_1951/type_cast_1937_Update/cr
      -- 
    rr_5158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(113), ack => type_cast_1937_inst_req_0); -- 
    cr_5163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(113), ack => type_cast_1937_inst_req_1); -- 
    zeropad3D_B_CP_4205_elements(113) <= OrReduce(zeropad3D_B_CP_4205_elements(50) & zeropad3D_B_CP_4205_elements(70));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	88 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Sample/$exit
      -- 
    ra_5608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	88 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/Update/$exit
      -- 
    ca_5613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	121 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_req
      -- CP-element group 116: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2066/$exit
      -- CP-element group 116: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2061/$exit
      -- 
    phi_stmt_2061_req_5614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2061_req_5614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(116), ack => phi_stmt_2061_req_1); -- 
    zeropad3D_B_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(114) & zeropad3D_B_CP_4205_elements(115);
      gj_zeropad3D_B_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  output  delay-element  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	88 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	121 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_req
      -- CP-element group 117: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2073_konst_delay_trans
      -- CP-element group 117: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2067/$exit
      -- 
    phi_stmt_2067_req_5622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2067_req_5622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(117), ack => phi_stmt_2067_req_1); -- 
    -- Element group zeropad3D_B_CP_4205_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_4205_elements(88), ack => zeropad3D_B_CP_4205_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Sample/$exit
      -- 
    ra_5639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2058_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	88 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Update/ca
      -- CP-element group 119: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/Update/$exit
      -- 
    ca_5644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2058_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/$exit
      -- CP-element group 120: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$exit
      -- CP-element group 120: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_req
      -- CP-element group 120: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/SplitProtocol/$exit
      -- CP-element group 120: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2058/$exit
      -- 
    phi_stmt_2055_req_5645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2055_req_5645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(120), ack => phi_stmt_2055_req_0); -- 
    zeropad3D_B_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(118) & zeropad3D_B_CP_4205_elements(119);
      gj_zeropad3D_B_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	116 
    -- CP-element group 121: 	117 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	132 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1483/ifx_xelse142_ifx_xend173_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(116) & zeropad3D_B_CP_4205_elements(117) & zeropad3D_B_CP_4205_elements(120);
      gj_zeropad3D_B_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	73 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/$exit
      -- 
    ra_5665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2064_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	73 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/ca
      -- CP-element group 123: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/$exit
      -- 
    ca_5670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2064_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	131 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_req
      -- CP-element group 124: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/$exit
      -- CP-element group 124: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/$exit
      -- CP-element group 124: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$exit
      -- CP-element group 124: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2061/$exit
      -- 
    phi_stmt_2061_req_5671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2061_req_5671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(124), ack => phi_stmt_2061_req_0); -- 
    zeropad3D_B_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(122) & zeropad3D_B_CP_4205_elements(123);
      gj_zeropad3D_B_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	73 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Sample/ra
      -- 
    ra_5688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2070_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	73 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Update/ca
      -- CP-element group 126: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/Update/$exit
      -- 
    ca_5693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2070_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	131 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/$exit
      -- CP-element group 127: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/$exit
      -- CP-element group 127: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/$exit
      -- CP-element group 127: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_sources/type_cast_2070/SplitProtocol/$exit
      -- CP-element group 127: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2067/phi_stmt_2067_req
      -- 
    phi_stmt_2067_req_5694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2067_req_5694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(127), ack => phi_stmt_2067_req_0); -- 
    zeropad3D_B_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(125) & zeropad3D_B_CP_4205_elements(126);
      gj_zeropad3D_B_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	73 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Sample/ra
      -- CP-element group 128: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Sample/$exit
      -- 
    ra_5711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2060_inst_ack_0, ack => zeropad3D_B_CP_4205_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	73 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Update/ca
      -- CP-element group 129: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/Update/$exit
      -- 
    ca_5716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2060_inst_ack_1, ack => zeropad3D_B_CP_4205_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_req
      -- CP-element group 130: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/SplitProtocol/$exit
      -- CP-element group 130: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/type_cast_2060/$exit
      -- CP-element group 130: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/phi_stmt_2055_sources/$exit
      -- CP-element group 130: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/phi_stmt_2055/$exit
      -- 
    phi_stmt_2055_req_5717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2055_req_5717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_4205_elements(130), ack => phi_stmt_2055_req_1); -- 
    zeropad3D_B_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(128) & zeropad3D_B_CP_4205_elements(129);
      gj_zeropad3D_B_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	124 
    -- CP-element group 131: 	127 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1483/ifx_xthen137_ifx_xend173_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(124) & zeropad3D_B_CP_4205_elements(127) & zeropad3D_B_CP_4205_elements(130);
      gj_zeropad3D_B_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  merge  fork  transition  place  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	121 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	135 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_1483/merge_stmt_2054_PhiAck/$entry
      -- CP-element group 132: 	 branch_block_stmt_1483/merge_stmt_2054_PhiReqMerge
      -- 
    zeropad3D_B_CP_4205_elements(132) <= OrReduce(zeropad3D_B_CP_4205_elements(121) & zeropad3D_B_CP_4205_elements(131));
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	136 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1483/merge_stmt_2054_PhiAck/phi_stmt_2055_ack
      -- 
    phi_stmt_2055_ack_5722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2055_ack_0, ack => zeropad3D_B_CP_4205_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1483/merge_stmt_2054_PhiAck/phi_stmt_2061_ack
      -- 
    phi_stmt_2061_ack_5723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2061_ack_0, ack => zeropad3D_B_CP_4205_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	132 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1483/merge_stmt_2054_PhiAck/phi_stmt_2067_ack
      -- 
    phi_stmt_2067_ack_5724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2067_ack_0, ack => zeropad3D_B_CP_4205_elements(135)); -- 
    -- CP-element group 136:  join  transition  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	133 
    -- CP-element group 136: 	134 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	1 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1483/merge_stmt_2054_PhiAck/$exit
      -- 
    zeropad3D_B_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_4205_elements(133) & zeropad3D_B_CP_4205_elements(134) & zeropad3D_B_CP_4205_elements(135);
      gj_zeropad3D_B_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_4205_elements(136), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1561_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1582_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1597_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1621_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1641_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1805_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1888_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1913_wire : std_logic_vector(31 downto 0);
    signal LOAD_pad_1511_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1511_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom122_1899_resized : std_logic_vector(13 downto 0);
    signal R_idxprom122_1899_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom127_1924_resized : std_logic_vector(13 downto 0);
    signal R_idxprom127_1924_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1816_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1816_scaled : std_logic_vector(13 downto 0);
    signal add103_1861 : std_logic_vector(31 downto 0);
    signal add113_1876 : std_logic_vector(31 downto 0);
    signal add119_1881 : std_logic_vector(31 downto 0);
    signal add132_1944 : std_logic_vector(31 downto 0);
    signal add140_1964 : std_logic_vector(15 downto 0);
    signal add149_1994 : std_logic_vector(31 downto 0);
    signal add164_2042 : std_logic_vector(31 downto 0);
    signal add65_1756 : std_logic_vector(31 downto 0);
    signal add76_1793 : std_logic_vector(31 downto 0);
    signal add82_1798 : std_logic_vector(31 downto 0);
    signal add94_1856 : std_logic_vector(31 downto 0);
    signal add_1708 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1817_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1817_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1817_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1817_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1817_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1817_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_root_address : std_logic_vector(13 downto 0);
    signal arrayidx123_1902 : std_logic_vector(31 downto 0);
    signal arrayidx128_1927 : std_logic_vector(31 downto 0);
    signal arrayidx_1819 : std_logic_vector(31 downto 0);
    signal call_1486 : std_logic_vector(15 downto 0);
    signal cmp135_1951 : std_logic_vector(0 downto 0);
    signal cmp150_1999 : std_logic_vector(0 downto 0);
    signal cmp165_2047 : std_logic_vector(0 downto 0);
    signal cmp50_1713 : std_logic_vector(0 downto 0);
    signal cmp57_1732 : std_logic_vector(0 downto 0);
    signal cmp66_1761 : std_logic_vector(0 downto 0);
    signal cmp_1678 : std_logic_vector(0 downto 0);
    signal conv131_1938 : std_logic_vector(31 downto 0);
    signal conv145_1977 : std_logic_vector(31 downto 0);
    signal conv158_2019 : std_logic_vector(31 downto 0);
    signal conv25_1563 : std_logic_vector(31 downto 0);
    signal conv31_1584 : std_logic_vector(31 downto 0);
    signal conv33_1599 : std_logic_vector(31 downto 0);
    signal conv40_1671 : std_logic_vector(31 downto 0);
    signal conv42_1608 : std_logic_vector(31 downto 0);
    signal conv54_1725 : std_logic_vector(31 downto 0);
    signal conv70_1773 : std_logic_vector(31 downto 0);
    signal conv74_1778 : std_logic_vector(31 downto 0);
    signal conv78_1623 : std_logic_vector(31 downto 0);
    signal conv86_1831 : std_logic_vector(31 downto 0);
    signal conv96_1643 : std_logic_vector(31 downto 0);
    signal conv_1509 : std_logic_vector(15 downto 0);
    signal div160_2037 : std_logic_vector(31 downto 0);
    signal div47_1703 : std_logic_vector(31 downto 0);
    signal div_1505 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1693 : std_logic_vector(31 downto 0);
    signal iNsTr_15_1985 : std_logic_vector(31 downto 0);
    signal iNsTr_16_2027 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1747 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1495 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1520 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1532 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1544 : std_logic_vector(31 downto 0);
    signal idxprom122_1895 : std_logic_vector(63 downto 0);
    signal idxprom127_1920 : std_logic_vector(63 downto 0);
    signal idxprom_1812 : std_logic_vector(63 downto 0);
    signal inc155_2003 : std_logic_vector(15 downto 0);
    signal inc155x_xix_x2_2008 : std_logic_vector(15 downto 0);
    signal inc_1972 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_2055 : std_logic_vector(15 downto 0);
    signal ix_x2_1646 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_2061 : std_logic_vector(15 downto 0);
    signal jx_x1_1653 : std_logic_vector(15 downto 0);
    signal jx_x2_2014 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_2067 : std_logic_vector(15 downto 0);
    signal kx_x1_1659 : std_logic_vector(15 downto 0);
    signal mul102_1851 : std_logic_vector(31 downto 0);
    signal mul112_1866 : std_logic_vector(31 downto 0);
    signal mul118_1871 : std_logic_vector(31 downto 0);
    signal mul34_1604 : std_logic_vector(31 downto 0);
    signal mul75_1783 : std_logic_vector(31 downto 0);
    signal mul81_1788 : std_logic_vector(31 downto 0);
    signal mul93_1841 : std_logic_vector(31 downto 0);
    signal ptr_deref_1498_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1498_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1498_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1498_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1498_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1523_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1535_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1535_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1535_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1535_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1535_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1547_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1547_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1547_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1547_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1547_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1696_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1696_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1696_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1696_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1696_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1750_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1750_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1750_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1750_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1750_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1821_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1821_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1821_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1821_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1821_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1821_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1905_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1929_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1929_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1929_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1929_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1929_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1929_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1988_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1988_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1988_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1988_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1988_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2030_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2030_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2030_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2030_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2030_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext175_1590 : std_logic_vector(31 downto 0);
    signal sext176_1634 : std_logic_vector(31 downto 0);
    signal sext182_1554 : std_logic_vector(31 downto 0);
    signal sext183_1575 : std_logic_vector(31 downto 0);
    signal sext184_1614 : std_logic_vector(31 downto 0);
    signal sext_1569 : std_logic_vector(31 downto 0);
    signal shl_1629 : std_logic_vector(31 downto 0);
    signal shr121_1890 : std_logic_vector(31 downto 0);
    signal shr126_1915 : std_logic_vector(31 downto 0);
    signal shr_1807 : std_logic_vector(31 downto 0);
    signal sub101_1846 : std_logic_vector(31 downto 0);
    signal sub_1836 : std_logic_vector(31 downto 0);
    signal tmp124_1906 : std_logic_vector(63 downto 0);
    signal tmp146_1989 : std_logic_vector(31 downto 0);
    signal tmp159_2031 : std_logic_vector(31 downto 0);
    signal tmp15_1536 : std_logic_vector(31 downto 0);
    signal tmp18_1548 : std_logic_vector(31 downto 0);
    signal tmp3_1512 : std_logic_vector(7 downto 0);
    signal tmp46_1697 : std_logic_vector(31 downto 0);
    signal tmp62_1751 : std_logic_vector(31 downto 0);
    signal tmp6_1524 : std_logic_vector(31 downto 0);
    signal tmp_1499 : std_logic_vector(31 downto 0);
    signal type_cast_1503_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1552_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1557_wire : std_logic_vector(31 downto 0);
    signal type_cast_1560_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1567_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1573_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1578_wire : std_logic_vector(31 downto 0);
    signal type_cast_1581_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1588_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1593_wire : std_logic_vector(31 downto 0);
    signal type_cast_1596_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1617_wire : std_logic_vector(31 downto 0);
    signal type_cast_1620_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1627_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1637_wire : std_logic_vector(31 downto 0);
    signal type_cast_1640_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1650_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1652_wire : std_logic_vector(15 downto 0);
    signal type_cast_1656_wire : std_logic_vector(15 downto 0);
    signal type_cast_1658_wire : std_logic_vector(15 downto 0);
    signal type_cast_1663_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1665_wire : std_logic_vector(15 downto 0);
    signal type_cast_1669_wire : std_logic_vector(31 downto 0);
    signal type_cast_1674_wire : std_logic_vector(31 downto 0);
    signal type_cast_1676_wire : std_logic_vector(31 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1723_wire : std_logic_vector(31 downto 0);
    signal type_cast_1728_wire : std_logic_vector(31 downto 0);
    signal type_cast_1730_wire : std_logic_vector(31 downto 0);
    signal type_cast_1771_wire : std_logic_vector(31 downto 0);
    signal type_cast_1776_wire : std_logic_vector(31 downto 0);
    signal type_cast_1801_wire : std_logic_vector(31 downto 0);
    signal type_cast_1804_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1810_wire : std_logic_vector(63 downto 0);
    signal type_cast_1823_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1829_wire : std_logic_vector(31 downto 0);
    signal type_cast_1884_wire : std_logic_vector(31 downto 0);
    signal type_cast_1887_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1893_wire : std_logic_vector(63 downto 0);
    signal type_cast_1909_wire : std_logic_vector(31 downto 0);
    signal type_cast_1912_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1918_wire : std_logic_vector(63 downto 0);
    signal type_cast_1936_wire : std_logic_vector(31 downto 0);
    signal type_cast_1942_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1947_wire : std_logic_vector(31 downto 0);
    signal type_cast_1949_wire : std_logic_vector(31 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1970_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1975_wire : std_logic_vector(31 downto 0);
    signal type_cast_2017_wire : std_logic_vector(31 downto 0);
    signal type_cast_2035_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2058_wire : std_logic_vector(15 downto 0);
    signal type_cast_2060_wire : std_logic_vector(15 downto 0);
    signal type_cast_2064_wire : std_logic_vector(15 downto 0);
    signal type_cast_2066_wire : std_logic_vector(15 downto 0);
    signal type_cast_2070_wire : std_logic_vector(15 downto 0);
    signal type_cast_2073_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_pad_1511_word_address_0 <= "0";
    array_obj_ref_1817_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1817_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1817_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1817_resized_base_address <= "00000000000000";
    array_obj_ref_1900_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1900_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1900_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1900_resized_base_address <= "00000000000000";
    array_obj_ref_1925_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1925_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1925_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1925_resized_base_address <= "00000000000000";
    iNsTr_10_1693 <= "00000000000000000000000000000011";
    iNsTr_15_1985 <= "00000000000000000000000000000100";
    iNsTr_16_2027 <= "00000000000000000000000000000011";
    iNsTr_18_1747 <= "00000000000000000000000000000100";
    iNsTr_2_1495 <= "00000000000000000000000000000100";
    iNsTr_3_1520 <= "00000000000000000000000000000101";
    iNsTr_4_1532 <= "00000000000000000000000000000101";
    iNsTr_5_1544 <= "00000000000000000000000000000100";
    ptr_deref_1498_word_offset_0 <= "0000000";
    ptr_deref_1523_word_offset_0 <= "0000000";
    ptr_deref_1535_word_offset_0 <= "0000000";
    ptr_deref_1547_word_offset_0 <= "0000000";
    ptr_deref_1696_word_offset_0 <= "0000000";
    ptr_deref_1750_word_offset_0 <= "0000000";
    ptr_deref_1821_word_offset_0 <= "00000000000000";
    ptr_deref_1905_word_offset_0 <= "00000000000000";
    ptr_deref_1929_word_offset_0 <= "00000000000000";
    ptr_deref_1988_word_offset_0 <= "0000000";
    ptr_deref_2030_word_offset_0 <= "0000000";
    type_cast_1503_wire_constant <= "00000000000000000000000000000001";
    type_cast_1552_wire_constant <= "00000000000000000000000000010000";
    type_cast_1560_wire_constant <= "00000000000000000000000000010000";
    type_cast_1567_wire_constant <= "00000000000000000000000000010000";
    type_cast_1573_wire_constant <= "00000000000000000000000000010000";
    type_cast_1581_wire_constant <= "00000000000000000000000000010000";
    type_cast_1588_wire_constant <= "00000000000000000000000000010000";
    type_cast_1596_wire_constant <= "00000000000000000000000000010000";
    type_cast_1612_wire_constant <= "00000000000000000000000000010000";
    type_cast_1620_wire_constant <= "00000000000000000000000000010000";
    type_cast_1627_wire_constant <= "00000000000000000000000000000001";
    type_cast_1640_wire_constant <= "00000000000000000000000000010000";
    type_cast_1650_wire_constant <= "0000000000000000";
    type_cast_1663_wire_constant <= "0000000000000000";
    type_cast_1701_wire_constant <= "00000000000000000000000000000001";
    type_cast_1804_wire_constant <= "00000000000000000000000000000010";
    type_cast_1823_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1887_wire_constant <= "00000000000000000000000000000010";
    type_cast_1912_wire_constant <= "00000000000000000000000000000010";
    type_cast_1942_wire_constant <= "00000000000000000000000000000100";
    type_cast_1962_wire_constant <= "0000000000000100";
    type_cast_1970_wire_constant <= "0000000000000001";
    type_cast_2035_wire_constant <= "00000000000000000000000000000001";
    type_cast_2073_wire_constant <= "0000000000000000";
    phi_stmt_1646: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1650_wire_constant & type_cast_1652_wire;
      req <= phi_stmt_1646_req_0 & phi_stmt_1646_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1646",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1646_ack_0,
          idata => idata,
          odata => ix_x2_1646,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1646
    phi_stmt_1653: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1656_wire & type_cast_1658_wire;
      req <= phi_stmt_1653_req_0 & phi_stmt_1653_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1653",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1653_ack_0,
          idata => idata,
          odata => jx_x1_1653,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1653
    phi_stmt_1659: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1663_wire_constant & type_cast_1665_wire;
      req <= phi_stmt_1659_req_0 & phi_stmt_1659_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1659",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1659_ack_0,
          idata => idata,
          odata => kx_x1_1659,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1659
    phi_stmt_2055: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2058_wire & type_cast_2060_wire;
      req <= phi_stmt_2055_req_0 & phi_stmt_2055_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2055",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2055_ack_0,
          idata => idata,
          odata => ix_x1x_xph_2055,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2055
    phi_stmt_2061: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2064_wire & type_cast_2066_wire;
      req <= phi_stmt_2061_req_0 & phi_stmt_2061_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2061",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2061_ack_0,
          idata => idata,
          odata => jx_x0x_xph_2061,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2061
    phi_stmt_2067: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2070_wire & type_cast_2073_wire_constant;
      req <= phi_stmt_2067_req_0 & phi_stmt_2067_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2067",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2067_ack_0,
          idata => idata,
          odata => kx_x0x_xph_2067,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2067
    -- flow-through select operator MUX_2013_inst
    jx_x2_2014 <= conv_1509 when (cmp150_1999(0) /=  '0') else inc_1972;
    addr_of_1818_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1818_final_reg_req_0;
      addr_of_1818_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1818_final_reg_req_1;
      addr_of_1818_final_reg_ack_1<= rack(0);
      addr_of_1818_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1818_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1817_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1819,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1901_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1901_final_reg_req_0;
      addr_of_1901_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1901_final_reg_req_1;
      addr_of_1901_final_reg_ack_1<= rack(0);
      addr_of_1901_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1901_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1900_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx123_1902,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1926_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1926_final_reg_req_0;
      addr_of_1926_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1926_final_reg_req_1;
      addr_of_1926_final_reg_ack_1<= rack(0);
      addr_of_1926_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1926_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1925_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx128_1927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1508_inst_req_0;
      type_cast_1508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1508_inst_req_1;
      type_cast_1508_inst_ack_1<= rack(0);
      type_cast_1508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1557_inst
    process(sext182_1554) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext182_1554(31 downto 0);
      type_cast_1557_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1562_inst
    process(ASHR_i32_i32_1561_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1561_wire(31 downto 0);
      conv25_1563 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1578_inst
    process(sext183_1575) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext183_1575(31 downto 0);
      type_cast_1578_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1583_inst
    process(ASHR_i32_i32_1582_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1582_wire(31 downto 0);
      conv31_1584 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1593_inst
    process(sext175_1590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext175_1590(31 downto 0);
      type_cast_1593_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1598_inst
    process(ASHR_i32_i32_1597_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1597_wire(31 downto 0);
      conv33_1599 <= tmp_var; -- 
    end process;
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1617_inst
    process(sext184_1614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext184_1614(31 downto 0);
      type_cast_1617_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1622_inst
    process(ASHR_i32_i32_1621_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1621_wire(31 downto 0);
      conv78_1623 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1637_inst
    process(sext176_1634) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext176_1634(31 downto 0);
      type_cast_1637_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1642_inst
    process(ASHR_i32_i32_1641_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1641_wire(31 downto 0);
      conv96_1643 <= tmp_var; -- 
    end process;
    type_cast_1652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1652_inst_req_0;
      type_cast_1652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1652_inst_req_1;
      type_cast_1652_inst_ack_1<= rack(0);
      type_cast_1652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_2055,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1652_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1656_inst_req_0;
      type_cast_1656_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1656_inst_req_1;
      type_cast_1656_inst_ack_1<= rack(0);
      type_cast_1656_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1656_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_1509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1656_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1658_inst_req_0;
      type_cast_1658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1658_inst_req_1;
      type_cast_1658_inst_ack_1<= rack(0);
      type_cast_1658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_2061,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1658_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1665_inst_req_0;
      type_cast_1665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1665_inst_req_1;
      type_cast_1665_inst_ack_1<= rack(0);
      type_cast_1665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_2067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1665_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1670_inst_req_0;
      type_cast_1670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1670_inst_req_1;
      type_cast_1670_inst_ack_1<= rack(0);
      type_cast_1670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1669_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_1671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1674_inst
    process(conv40_1671) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv40_1671(31 downto 0);
      type_cast_1674_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1676_inst
    process(conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv42_1608(31 downto 0);
      type_cast_1676_wire <= tmp_var; -- 
    end process;
    type_cast_1724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1724_inst_req_0;
      type_cast_1724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1724_inst_req_1;
      type_cast_1724_inst_ack_1<= rack(0);
      type_cast_1724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1723_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_1725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1728_inst
    process(conv54_1725) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv54_1725(31 downto 0);
      type_cast_1728_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1730_inst
    process(conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv42_1608(31 downto 0);
      type_cast_1730_wire <= tmp_var; -- 
    end process;
    type_cast_1772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1772_inst_req_0;
      type_cast_1772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1772_inst_req_1;
      type_cast_1772_inst_ack_1<= rack(0);
      type_cast_1772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1771_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1777_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1777_inst_req_0;
      type_cast_1777_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1777_inst_req_1;
      type_cast_1777_inst_ack_1<= rack(0);
      type_cast_1777_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1777_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1776_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1778,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1801_inst
    process(add82_1798) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add82_1798(31 downto 0);
      type_cast_1801_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1806_inst
    process(ASHR_i32_i32_1805_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1805_wire(31 downto 0);
      shr_1807 <= tmp_var; -- 
    end process;
    type_cast_1811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1811_inst_req_0;
      type_cast_1811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1811_inst_req_1;
      type_cast_1811_inst_ack_1<= rack(0);
      type_cast_1811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1810_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1812,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1830_inst_req_0;
      type_cast_1830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1830_inst_req_1;
      type_cast_1830_inst_ack_1<= rack(0);
      type_cast_1830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1829_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_1831,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1884_inst
    process(add103_1861) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add103_1861(31 downto 0);
      type_cast_1884_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1889_inst
    process(ASHR_i32_i32_1888_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1888_wire(31 downto 0);
      shr121_1890 <= tmp_var; -- 
    end process;
    type_cast_1894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1894_inst_req_0;
      type_cast_1894_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1894_inst_req_1;
      type_cast_1894_inst_ack_1<= rack(0);
      type_cast_1894_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1894_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1893_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom122_1895,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1909_inst
    process(add119_1881) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add119_1881(31 downto 0);
      type_cast_1909_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1914_inst
    process(ASHR_i32_i32_1913_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1913_wire(31 downto 0);
      shr126_1915 <= tmp_var; -- 
    end process;
    type_cast_1919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1919_inst_req_0;
      type_cast_1919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1919_inst_req_1;
      type_cast_1919_inst_ack_1<= rack(0);
      type_cast_1919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1918_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom127_1920,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1937_inst_req_0;
      type_cast_1937_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1937_inst_req_1;
      type_cast_1937_inst_ack_1<= rack(0);
      type_cast_1937_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1937_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1936_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_1938,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1947_inst
    process(add132_1944) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add132_1944(31 downto 0);
      type_cast_1947_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1949_inst
    process(conv25_1563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv25_1563(31 downto 0);
      type_cast_1949_wire <= tmp_var; -- 
    end process;
    type_cast_1976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1976_inst_req_0;
      type_cast_1976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1976_inst_req_1;
      type_cast_1976_inst_ack_1<= rack(0);
      type_cast_1976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1975_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2002_inst_req_0;
      type_cast_2002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2002_inst_req_1;
      type_cast_2002_inst_ack_1<= rack(0);
      type_cast_2002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2002_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp150_1999,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc155_2003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2018_inst_req_0;
      type_cast_2018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2018_inst_req_1;
      type_cast_2018_inst_ack_1<= rack(0);
      type_cast_2018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2017_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_2019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2058_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2058_inst_req_0;
      type_cast_2058_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2058_inst_req_1;
      type_cast_2058_inst_ack_1<= rack(0);
      type_cast_2058_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2058_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc155x_xix_x2_2008,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2058_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2060_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2060_inst_req_0;
      type_cast_2060_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2060_inst_req_1;
      type_cast_2060_inst_ack_1<= rack(0);
      type_cast_2060_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2060_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_1646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2060_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2064_inst_req_0;
      type_cast_2064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2064_inst_req_1;
      type_cast_2064_inst_ack_1<= rack(0);
      type_cast_2064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_1653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2064_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2066_inst_req_0;
      type_cast_2066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2066_inst_req_1;
      type_cast_2066_inst_ack_1<= rack(0);
      type_cast_2066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_2014,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2066_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2070_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2070_inst_req_0;
      type_cast_2070_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2070_inst_req_1;
      type_cast_2070_inst_ack_1<= rack(0);
      type_cast_2070_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2070_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add140_1964,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2070_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_pad_1511_gather_scatter
    process(LOAD_pad_1511_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1511_data_0;
      ov(7 downto 0) := iv;
      tmp3_1512 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1817_index_1_rename
    process(R_idxprom_1816_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1816_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1816_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1817_index_1_resize
    process(idxprom_1812) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1812;
      ov := iv(13 downto 0);
      R_idxprom_1816_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1817_root_address_inst
    process(array_obj_ref_1817_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1817_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1817_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1900_index_1_rename
    process(R_idxprom122_1899_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom122_1899_resized;
      ov(13 downto 0) := iv;
      R_idxprom122_1899_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1900_index_1_resize
    process(idxprom122_1895) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom122_1895;
      ov := iv(13 downto 0);
      R_idxprom122_1899_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1900_root_address_inst
    process(array_obj_ref_1900_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1900_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1900_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1925_index_1_rename
    process(R_idxprom127_1924_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom127_1924_resized;
      ov(13 downto 0) := iv;
      R_idxprom127_1924_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1925_index_1_resize
    process(idxprom127_1920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom127_1920;
      ov := iv(13 downto 0);
      R_idxprom127_1924_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1925_root_address_inst
    process(array_obj_ref_1925_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1925_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1925_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1498_addr_0
    process(ptr_deref_1498_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1498_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1498_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1498_base_resize
    process(iNsTr_2_1495) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1495;
      ov := iv(6 downto 0);
      ptr_deref_1498_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1498_gather_scatter
    process(ptr_deref_1498_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1498_data_0;
      ov(31 downto 0) := iv;
      tmp_1499 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1498_root_address_inst
    process(ptr_deref_1498_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1498_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1498_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_addr_0
    process(ptr_deref_1523_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1523_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1523_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_base_resize
    process(iNsTr_3_1520) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1520;
      ov := iv(6 downto 0);
      ptr_deref_1523_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_gather_scatter
    process(ptr_deref_1523_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1523_data_0;
      ov(31 downto 0) := iv;
      tmp6_1524 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_root_address_inst
    process(ptr_deref_1523_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1523_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1523_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_addr_0
    process(ptr_deref_1535_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1535_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1535_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_base_resize
    process(iNsTr_4_1532) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1532;
      ov := iv(6 downto 0);
      ptr_deref_1535_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_gather_scatter
    process(ptr_deref_1535_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1535_data_0;
      ov(31 downto 0) := iv;
      tmp15_1536 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1535_root_address_inst
    process(ptr_deref_1535_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1535_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1535_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_addr_0
    process(ptr_deref_1547_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1547_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1547_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_base_resize
    process(iNsTr_5_1544) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1544;
      ov := iv(6 downto 0);
      ptr_deref_1547_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_gather_scatter
    process(ptr_deref_1547_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1547_data_0;
      ov(31 downto 0) := iv;
      tmp18_1548 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1547_root_address_inst
    process(ptr_deref_1547_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1547_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1547_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1696_addr_0
    process(ptr_deref_1696_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1696_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1696_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1696_base_resize
    process(iNsTr_10_1693) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1693;
      ov := iv(6 downto 0);
      ptr_deref_1696_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1696_gather_scatter
    process(ptr_deref_1696_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1696_data_0;
      ov(31 downto 0) := iv;
      tmp46_1697 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1696_root_address_inst
    process(ptr_deref_1696_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1696_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1696_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_addr_0
    process(ptr_deref_1750_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1750_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1750_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_base_resize
    process(iNsTr_18_1747) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_1747;
      ov := iv(6 downto 0);
      ptr_deref_1750_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_gather_scatter
    process(ptr_deref_1750_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1750_data_0;
      ov(31 downto 0) := iv;
      tmp62_1751 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_root_address_inst
    process(ptr_deref_1750_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1750_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1750_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1821_addr_0
    process(ptr_deref_1821_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1821_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1821_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1821_base_resize
    process(arrayidx_1819) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1819;
      ov := iv(13 downto 0);
      ptr_deref_1821_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1821_gather_scatter
    process(type_cast_1823_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1823_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1821_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1821_root_address_inst
    process(ptr_deref_1821_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1821_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1821_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_addr_0
    process(ptr_deref_1905_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1905_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_base_resize
    process(arrayidx123_1902) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx123_1902;
      ov := iv(13 downto 0);
      ptr_deref_1905_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_gather_scatter
    process(ptr_deref_1905_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_data_0;
      ov(63 downto 0) := iv;
      tmp124_1906 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_root_address_inst
    process(ptr_deref_1905_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1905_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1929_addr_0
    process(ptr_deref_1929_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1929_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1929_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1929_base_resize
    process(arrayidx128_1927) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx128_1927;
      ov := iv(13 downto 0);
      ptr_deref_1929_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1929_gather_scatter
    process(tmp124_1906) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp124_1906;
      ov(63 downto 0) := iv;
      ptr_deref_1929_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1929_root_address_inst
    process(ptr_deref_1929_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1929_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1929_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1988_addr_0
    process(ptr_deref_1988_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1988_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1988_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1988_base_resize
    process(iNsTr_15_1985) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_1985;
      ov := iv(6 downto 0);
      ptr_deref_1988_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1988_gather_scatter
    process(ptr_deref_1988_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1988_data_0;
      ov(31 downto 0) := iv;
      tmp146_1989 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1988_root_address_inst
    process(ptr_deref_1988_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1988_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1988_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2030_addr_0
    process(ptr_deref_2030_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2030_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2030_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2030_base_resize
    process(iNsTr_16_2027) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_16_2027;
      ov := iv(6 downto 0);
      ptr_deref_2030_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2030_gather_scatter
    process(ptr_deref_2030_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2030_data_0;
      ov(31 downto 0) := iv;
      tmp159_2031 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2030_root_address_inst
    process(ptr_deref_2030_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2030_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2030_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1679_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1678;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1679_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1679_branch_req_0,
          ack0 => if_stmt_1679_branch_ack_0,
          ack1 => if_stmt_1679_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1714_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp50_1713;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1714_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1714_branch_req_0,
          ack0 => if_stmt_1714_branch_ack_0,
          ack1 => if_stmt_1714_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1733_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp57_1732;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1733_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1733_branch_req_0,
          ack0 => if_stmt_1733_branch_ack_0,
          ack1 => if_stmt_1733_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1762_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp66_1761;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1762_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1762_branch_req_0,
          ack0 => if_stmt_1762_branch_ack_0,
          ack1 => if_stmt_1762_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1952_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp135_1951;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1952_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1952_branch_req_0,
          ack0 => if_stmt_1952_branch_ack_0,
          ack1 => if_stmt_1952_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2048_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp165_2047;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2048_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2048_branch_req_0,
          ack0 => if_stmt_2048_branch_ack_0,
          ack1 => if_stmt_2048_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1963_inst
    process(kx_x1_1659) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_1659, type_cast_1962_wire_constant, tmp_var);
      add140_1964 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1971_inst
    process(jx_x1_1653) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_1653, type_cast_1970_wire_constant, tmp_var);
      inc_1972 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2007_inst
    process(inc155_2003, ix_x2_1646) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc155_2003, ix_x2_1646, tmp_var);
      inc155x_xix_x2_2008 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1707_inst
    process(div47_1703, conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div47_1703, conv42_1608, tmp_var);
      add_1708 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1755_inst
    process(tmp62_1751, conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp62_1751, conv42_1608, tmp_var);
      add65_1756 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1792_inst
    process(mul75_1783, mul81_1788) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul75_1783, mul81_1788, tmp_var);
      add76_1793 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1797_inst
    process(add76_1793, conv70_1773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add76_1793, conv70_1773, tmp_var);
      add82_1798 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1855_inst
    process(conv86_1831, mul102_1851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv86_1831, mul102_1851, tmp_var);
      add94_1856 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1860_inst
    process(add94_1856, mul93_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add94_1856, mul93_1841, tmp_var);
      add103_1861 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1875_inst
    process(mul112_1866, mul118_1871) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul112_1866, mul118_1871, tmp_var);
      add113_1876 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1880_inst
    process(add113_1876, conv86_1831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add113_1876, conv86_1831, tmp_var);
      add119_1881 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1943_inst
    process(conv131_1938) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv131_1938, type_cast_1942_wire_constant, tmp_var);
      add132_1944 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1993_inst
    process(tmp146_1989, shl_1629) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp146_1989, shl_1629, tmp_var);
      add149_1994 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2041_inst
    process(div160_2037, shl_1629) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div160_2037, shl_1629, tmp_var);
      add164_2042 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1561_inst
    process(type_cast_1557_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1557_wire, type_cast_1560_wire_constant, tmp_var);
      ASHR_i32_i32_1561_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1582_inst
    process(type_cast_1578_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1578_wire, type_cast_1581_wire_constant, tmp_var);
      ASHR_i32_i32_1582_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1597_inst
    process(type_cast_1593_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1593_wire, type_cast_1596_wire_constant, tmp_var);
      ASHR_i32_i32_1597_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1621_inst
    process(type_cast_1617_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1617_wire, type_cast_1620_wire_constant, tmp_var);
      ASHR_i32_i32_1621_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1641_inst
    process(type_cast_1637_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1637_wire, type_cast_1640_wire_constant, tmp_var);
      ASHR_i32_i32_1641_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1805_inst
    process(type_cast_1801_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1801_wire, type_cast_1804_wire_constant, tmp_var);
      ASHR_i32_i32_1805_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1888_inst
    process(type_cast_1884_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1884_wire, type_cast_1887_wire_constant, tmp_var);
      ASHR_i32_i32_1888_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1913_inst
    process(type_cast_1909_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1909_wire, type_cast_1912_wire_constant, tmp_var);
      ASHR_i32_i32_1913_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1998_inst
    process(conv145_1977, add149_1994) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv145_1977, add149_1994, tmp_var);
      cmp150_1999 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2046_inst
    process(conv158_2019, add164_2042) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv158_2019, add164_2042, tmp_var);
      cmp165_2047 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1504_inst
    process(tmp_1499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1499, type_cast_1503_wire_constant, tmp_var);
      div_1505 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1702_inst
    process(tmp46_1697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp46_1697, type_cast_1701_wire_constant, tmp_var);
      div47_1703 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2036_inst
    process(tmp159_2031) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp159_2031, type_cast_2035_wire_constant, tmp_var);
      div160_2037 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1603_inst
    process(conv33_1599, conv31_1584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_1599, conv31_1584, tmp_var);
      mul34_1604 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1633_inst
    process(sext_1569, conv25_1563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sext_1569, conv25_1563, tmp_var);
      sext176_1634 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1782_inst
    process(conv74_1778, conv31_1584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv74_1778, conv31_1584, tmp_var);
      mul75_1783 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1787_inst
    process(conv40_1671, conv78_1623) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv40_1671, conv78_1623, tmp_var);
      mul81_1788 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1840_inst
    process(sub_1836, conv25_1563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1836, conv25_1563, tmp_var);
      mul93_1841 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1850_inst
    process(sub101_1846, conv96_1643) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub101_1846, conv96_1643, tmp_var);
      mul102_1851 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1865_inst
    process(conv54_1725, conv31_1584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv54_1725, conv31_1584, tmp_var);
      mul112_1866 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1870_inst
    process(conv40_1671, conv78_1623) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv40_1671, conv78_1623, tmp_var);
      mul118_1871 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1553_inst
    process(tmp6_1524) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp6_1524, type_cast_1552_wire_constant, tmp_var);
      sext182_1554 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1568_inst
    process(tmp_1499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp_1499, type_cast_1567_wire_constant, tmp_var);
      sext_1569 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1574_inst
    process(tmp15_1536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp15_1536, type_cast_1573_wire_constant, tmp_var);
      sext183_1575 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1589_inst
    process(tmp18_1548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp18_1548, type_cast_1588_wire_constant, tmp_var);
      sext175_1590 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1613_inst
    process(mul34_1604) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul34_1604, type_cast_1612_wire_constant, tmp_var);
      sext184_1614 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1628_inst
    process(conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv42_1608, type_cast_1627_wire_constant, tmp_var);
      shl_1629 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1677_inst
    process(type_cast_1674_wire, type_cast_1676_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1674_wire, type_cast_1676_wire, tmp_var);
      cmp_1678 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1731_inst
    process(type_cast_1728_wire, type_cast_1730_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1728_wire, type_cast_1730_wire, tmp_var);
      cmp57_1732 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1950_inst
    process(type_cast_1947_wire, type_cast_1949_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1947_wire, type_cast_1949_wire, tmp_var);
      cmp135_1951 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1835_inst
    process(conv54_1725, conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv54_1725, conv42_1608, tmp_var);
      sub_1836 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1845_inst
    process(conv40_1671, conv42_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv40_1671, conv42_1608, tmp_var);
      sub101_1846 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1712_inst
    process(conv40_1671, add_1708) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv40_1671, add_1708, tmp_var);
      cmp50_1713 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1760_inst
    process(conv54_1725, add65_1756) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv54_1725, add65_1756, tmp_var);
      cmp66_1761 <= tmp_var; --
    end process;
    -- shared split operator group (48) : array_obj_ref_1817_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1816_scaled;
      array_obj_ref_1817_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1817_index_offset_req_0;
      array_obj_ref_1817_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1817_index_offset_req_1;
      array_obj_ref_1817_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : array_obj_ref_1900_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom122_1899_scaled;
      array_obj_ref_1900_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1900_index_offset_req_0;
      array_obj_ref_1900_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1900_index_offset_req_1;
      array_obj_ref_1900_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : array_obj_ref_1925_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom127_1924_scaled;
      array_obj_ref_1925_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1925_index_offset_req_0;
      array_obj_ref_1925_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1925_index_offset_req_1;
      array_obj_ref_1925_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- unary operator type_cast_1669_inst
    process(ix_x2_1646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_1646, tmp_var);
      type_cast_1669_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1723_inst
    process(jx_x1_1653) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1653, tmp_var);
      type_cast_1723_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1771_inst
    process(kx_x1_1659) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1659, tmp_var);
      type_cast_1771_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1776_inst
    process(jx_x1_1653) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1653, tmp_var);
      type_cast_1776_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1810_inst
    process(shr_1807) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1807, tmp_var);
      type_cast_1810_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1829_inst
    process(kx_x1_1659) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1659, tmp_var);
      type_cast_1829_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1893_inst
    process(shr121_1890) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr121_1890, tmp_var);
      type_cast_1893_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1918_inst
    process(shr126_1915) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr126_1915, tmp_var);
      type_cast_1918_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1936_inst
    process(kx_x1_1659) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1659, tmp_var);
      type_cast_1936_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1975_inst
    process(inc_1972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1972, tmp_var);
      type_cast_1975_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2017_inst
    process(inc155x_xix_x2_2008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc155x_xix_x2_2008, tmp_var);
      type_cast_2017_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_pad_1511_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_pad_1511_load_0_req_0;
      LOAD_pad_1511_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_pad_1511_load_0_req_1;
      LOAD_pad_1511_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_1511_word_address_0;
      LOAD_pad_1511_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(0 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1750_load_0 ptr_deref_1988_load_0 ptr_deref_2030_load_0 ptr_deref_1696_load_0 ptr_deref_1498_load_0 ptr_deref_1523_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(41 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_1750_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1988_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2030_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1696_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1498_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1523_load_0_req_0;
      ptr_deref_1750_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1988_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2030_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1696_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1498_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1523_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_1750_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1988_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2030_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1696_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1498_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1523_load_0_req_1;
      ptr_deref_1750_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1988_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2030_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1696_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1498_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1523_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1750_word_address_0 & ptr_deref_1988_word_address_0 & ptr_deref_2030_word_address_0 & ptr_deref_1696_word_address_0 & ptr_deref_1498_word_address_0 & ptr_deref_1523_word_address_0;
      ptr_deref_1750_data_0 <= data_out(191 downto 160);
      ptr_deref_1988_data_0 <= data_out(159 downto 128);
      ptr_deref_2030_data_0 <= data_out(127 downto 96);
      ptr_deref_1696_data_0 <= data_out(95 downto 64);
      ptr_deref_1498_data_0 <= data_out(63 downto 32);
      ptr_deref_1523_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1535_load_0 ptr_deref_1547_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1535_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1547_load_0_req_0;
      ptr_deref_1535_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1547_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1535_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1547_load_0_req_1;
      ptr_deref_1535_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1547_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1535_word_address_0 & ptr_deref_1547_word_address_0;
      ptr_deref_1535_data_0 <= data_out(63 downto 32);
      ptr_deref_1547_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(6 downto 0),
          mtag => memory_space_4_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1905_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1905_load_0_req_0;
      ptr_deref_1905_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1905_load_0_req_1;
      ptr_deref_1905_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1905_word_address_0;
      ptr_deref_1905_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_1821_store_0 ptr_deref_1929_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1821_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1929_store_0_req_0;
      ptr_deref_1821_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1929_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1821_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1929_store_0_req_1;
      ptr_deref_1821_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1929_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1821_word_address_0 & ptr_deref_1929_word_address_0;
      data_in <= ptr_deref_1821_data_0 & ptr_deref_1929_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_starting_1485_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_starting_1485_inst_req_0;
      RPIPE_Block1_starting_1485_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_starting_1485_inst_req_1;
      RPIPE_Block1_starting_1485_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1486 <= data_out(15 downto 0);
      Block1_starting_read_0_gI: SplitGuardInterface generic map(name => "Block1_starting_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block1_starting_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_starting_pipe_read_req(0),
          oack => Block1_starting_pipe_read_ack(0),
          odata => Block1_starting_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_complete_2078_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_complete_2078_inst_req_0;
      WPIPE_Block1_complete_2078_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_complete_2078_inst_req_1;
      WPIPE_Block1_complete_2078_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1486;
      Block1_complete_write_0_gI: SplitGuardInterface generic map(name => "Block1_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_complete", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_complete_pipe_write_req(0),
          oack => Block1_complete_pipe_write_ack(0),
          odata => Block1_complete_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_B_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_C is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block2_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_C;
architecture zeropad3D_C_arch of zeropad3D_C is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_C_CP_5741_start: Boolean;
  signal zeropad3D_C_CP_5741_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2138_load_0_ack_0 : boolean;
  signal type_cast_2111_inst_req_0 : boolean;
  signal ptr_deref_2126_load_0_req_1 : boolean;
  signal ptr_deref_2126_load_0_ack_1 : boolean;
  signal type_cast_2111_inst_ack_0 : boolean;
  signal ptr_deref_2138_load_0_req_0 : boolean;
  signal ptr_deref_2126_load_0_req_0 : boolean;
  signal ptr_deref_2126_load_0_ack_0 : boolean;
  signal ptr_deref_2138_load_0_req_1 : boolean;
  signal ptr_deref_2138_load_0_ack_1 : boolean;
  signal ptr_deref_2150_load_0_ack_0 : boolean;
  signal type_cast_2295_inst_ack_0 : boolean;
  signal phi_stmt_2692_req_0 : boolean;
  signal type_cast_2111_inst_req_1 : boolean;
  signal type_cast_2111_inst_ack_1 : boolean;
  signal ptr_deref_2150_load_0_req_0 : boolean;
  signal LOAD_pad_2114_load_0_req_0 : boolean;
  signal ptr_deref_2101_load_0_req_0 : boolean;
  signal ptr_deref_2101_load_0_ack_0 : boolean;
  signal LOAD_pad_2114_load_0_ack_0 : boolean;
  signal ptr_deref_2150_load_0_req_1 : boolean;
  signal ptr_deref_2150_load_0_ack_1 : boolean;
  signal phi_stmt_2282_req_1 : boolean;
  signal LOAD_pad_2114_load_0_ack_1 : boolean;
  signal type_cast_2697_inst_ack_0 : boolean;
  signal ptr_deref_2101_load_0_ack_1 : boolean;
  signal LOAD_pad_2114_load_0_req_1 : boolean;
  signal ptr_deref_2162_load_0_req_0 : boolean;
  signal ptr_deref_2162_load_0_ack_0 : boolean;
  signal type_cast_2295_inst_req_0 : boolean;
  signal ptr_deref_2101_load_0_req_1 : boolean;
  signal type_cast_2295_inst_req_1 : boolean;
  signal type_cast_2295_inst_ack_1 : boolean;
  signal type_cast_2697_inst_req_1 : boolean;
  signal type_cast_2697_inst_ack_1 : boolean;
  signal type_cast_2701_inst_req_0 : boolean;
  signal type_cast_2689_inst_req_0 : boolean;
  signal type_cast_2689_inst_ack_0 : boolean;
  signal phi_stmt_2692_req_1 : boolean;
  signal RPIPE_Block2_starting_2088_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_2088_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_2088_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_2088_inst_ack_1 : boolean;
  signal ptr_deref_2162_load_0_req_1 : boolean;
  signal ptr_deref_2162_load_0_ack_1 : boolean;
  signal type_cast_2216_inst_req_0 : boolean;
  signal type_cast_2216_inst_ack_0 : boolean;
  signal type_cast_2216_inst_req_1 : boolean;
  signal type_cast_2216_inst_ack_1 : boolean;
  signal type_cast_2300_inst_req_0 : boolean;
  signal type_cast_2300_inst_ack_0 : boolean;
  signal type_cast_2300_inst_req_1 : boolean;
  signal type_cast_2300_inst_ack_1 : boolean;
  signal if_stmt_2309_branch_req_0 : boolean;
  signal if_stmt_2309_branch_ack_1 : boolean;
  signal if_stmt_2309_branch_ack_0 : boolean;
  signal ptr_deref_2326_load_0_req_0 : boolean;
  signal ptr_deref_2326_load_0_ack_0 : boolean;
  signal ptr_deref_2326_load_0_req_1 : boolean;
  signal ptr_deref_2326_load_0_ack_1 : boolean;
  signal if_stmt_2338_branch_req_0 : boolean;
  signal if_stmt_2338_branch_ack_1 : boolean;
  signal if_stmt_2338_branch_ack_0 : boolean;
  signal type_cast_2348_inst_req_0 : boolean;
  signal type_cast_2348_inst_ack_0 : boolean;
  signal type_cast_2348_inst_req_1 : boolean;
  signal type_cast_2348_inst_ack_1 : boolean;
  signal if_stmt_2357_branch_req_0 : boolean;
  signal if_stmt_2357_branch_ack_1 : boolean;
  signal if_stmt_2357_branch_ack_0 : boolean;
  signal ptr_deref_2374_load_0_req_0 : boolean;
  signal ptr_deref_2374_load_0_ack_0 : boolean;
  signal ptr_deref_2374_load_0_req_1 : boolean;
  signal ptr_deref_2374_load_0_ack_1 : boolean;
  signal if_stmt_2392_branch_req_0 : boolean;
  signal if_stmt_2392_branch_ack_1 : boolean;
  signal if_stmt_2392_branch_ack_0 : boolean;
  signal type_cast_2402_inst_req_0 : boolean;
  signal type_cast_2402_inst_ack_0 : boolean;
  signal type_cast_2402_inst_req_1 : boolean;
  signal type_cast_2402_inst_ack_1 : boolean;
  signal type_cast_2407_inst_req_0 : boolean;
  signal type_cast_2407_inst_ack_0 : boolean;
  signal type_cast_2407_inst_req_1 : boolean;
  signal type_cast_2407_inst_ack_1 : boolean;
  signal type_cast_2441_inst_req_0 : boolean;
  signal type_cast_2441_inst_ack_0 : boolean;
  signal type_cast_2441_inst_req_1 : boolean;
  signal type_cast_2441_inst_ack_1 : boolean;
  signal phi_stmt_2686_req_0 : boolean;
  signal type_cast_2288_inst_ack_1 : boolean;
  signal type_cast_2697_inst_req_0 : boolean;
  signal array_obj_ref_2447_index_offset_req_0 : boolean;
  signal array_obj_ref_2447_index_offset_ack_0 : boolean;
  signal array_obj_ref_2447_index_offset_req_1 : boolean;
  signal array_obj_ref_2447_index_offset_ack_1 : boolean;
  signal type_cast_2695_inst_ack_1 : boolean;
  signal addr_of_2448_final_reg_req_0 : boolean;
  signal addr_of_2448_final_reg_ack_0 : boolean;
  signal type_cast_2288_inst_req_1 : boolean;
  signal type_cast_2695_inst_req_1 : boolean;
  signal addr_of_2448_final_reg_req_1 : boolean;
  signal phi_stmt_2686_req_1 : boolean;
  signal addr_of_2448_final_reg_ack_1 : boolean;
  signal type_cast_2689_inst_ack_1 : boolean;
  signal type_cast_2689_inst_req_1 : boolean;
  signal type_cast_2691_inst_ack_1 : boolean;
  signal type_cast_2691_inst_req_1 : boolean;
  signal ptr_deref_2451_store_0_req_0 : boolean;
  signal ptr_deref_2451_store_0_ack_0 : boolean;
  signal ptr_deref_2451_store_0_req_1 : boolean;
  signal ptr_deref_2451_store_0_ack_1 : boolean;
  signal type_cast_2691_inst_ack_0 : boolean;
  signal phi_stmt_2289_ack_0 : boolean;
  signal phi_stmt_2282_ack_0 : boolean;
  signal type_cast_2288_inst_ack_0 : boolean;
  signal type_cast_2691_inst_req_0 : boolean;
  signal type_cast_2460_inst_req_0 : boolean;
  signal type_cast_2460_inst_ack_0 : boolean;
  signal type_cast_2695_inst_ack_0 : boolean;
  signal type_cast_2460_inst_req_1 : boolean;
  signal type_cast_2460_inst_ack_1 : boolean;
  signal phi_stmt_2276_ack_0 : boolean;
  signal type_cast_2695_inst_req_0 : boolean;
  signal type_cast_2524_inst_req_0 : boolean;
  signal type_cast_2524_inst_ack_0 : boolean;
  signal type_cast_2288_inst_req_0 : boolean;
  signal type_cast_2524_inst_req_1 : boolean;
  signal type_cast_2524_inst_ack_1 : boolean;
  signal phi_stmt_2289_req_1 : boolean;
  signal phi_stmt_2698_req_1 : boolean;
  signal array_obj_ref_2530_index_offset_req_0 : boolean;
  signal array_obj_ref_2530_index_offset_ack_0 : boolean;
  signal array_obj_ref_2530_index_offset_req_1 : boolean;
  signal array_obj_ref_2530_index_offset_ack_1 : boolean;
  signal addr_of_2531_final_reg_req_0 : boolean;
  signal addr_of_2531_final_reg_ack_0 : boolean;
  signal addr_of_2531_final_reg_req_1 : boolean;
  signal addr_of_2531_final_reg_ack_1 : boolean;
  signal ptr_deref_2535_load_0_req_0 : boolean;
  signal ptr_deref_2535_load_0_ack_0 : boolean;
  signal ptr_deref_2535_load_0_req_1 : boolean;
  signal ptr_deref_2535_load_0_ack_1 : boolean;
  signal type_cast_2549_inst_req_0 : boolean;
  signal type_cast_2549_inst_ack_0 : boolean;
  signal type_cast_2549_inst_req_1 : boolean;
  signal type_cast_2549_inst_ack_1 : boolean;
  signal array_obj_ref_2555_index_offset_req_0 : boolean;
  signal array_obj_ref_2555_index_offset_ack_0 : boolean;
  signal array_obj_ref_2555_index_offset_req_1 : boolean;
  signal array_obj_ref_2555_index_offset_ack_1 : boolean;
  signal addr_of_2556_final_reg_req_0 : boolean;
  signal addr_of_2556_final_reg_ack_0 : boolean;
  signal addr_of_2556_final_reg_req_1 : boolean;
  signal addr_of_2556_final_reg_ack_1 : boolean;
  signal ptr_deref_2559_store_0_req_0 : boolean;
  signal ptr_deref_2559_store_0_ack_0 : boolean;
  signal ptr_deref_2559_store_0_req_1 : boolean;
  signal ptr_deref_2559_store_0_ack_1 : boolean;
  signal type_cast_2567_inst_req_0 : boolean;
  signal type_cast_2567_inst_ack_0 : boolean;
  signal type_cast_2567_inst_req_1 : boolean;
  signal type_cast_2567_inst_ack_1 : boolean;
  signal if_stmt_2582_branch_req_0 : boolean;
  signal if_stmt_2582_branch_ack_1 : boolean;
  signal if_stmt_2582_branch_ack_0 : boolean;
  signal type_cast_2606_inst_req_0 : boolean;
  signal type_cast_2606_inst_ack_0 : boolean;
  signal type_cast_2606_inst_req_1 : boolean;
  signal type_cast_2606_inst_ack_1 : boolean;
  signal ptr_deref_2618_load_0_req_0 : boolean;
  signal ptr_deref_2618_load_0_ack_0 : boolean;
  signal ptr_deref_2618_load_0_req_1 : boolean;
  signal ptr_deref_2618_load_0_ack_1 : boolean;
  signal type_cast_2638_inst_req_0 : boolean;
  signal type_cast_2638_inst_ack_0 : boolean;
  signal type_cast_2638_inst_req_1 : boolean;
  signal type_cast_2638_inst_ack_1 : boolean;
  signal type_cast_2655_inst_req_0 : boolean;
  signal type_cast_2655_inst_ack_0 : boolean;
  signal type_cast_2655_inst_req_1 : boolean;
  signal type_cast_2655_inst_ack_1 : boolean;
  signal ptr_deref_2667_load_0_req_0 : boolean;
  signal ptr_deref_2667_load_0_ack_0 : boolean;
  signal ptr_deref_2667_load_0_req_1 : boolean;
  signal ptr_deref_2667_load_0_ack_1 : boolean;
  signal if_stmt_2679_branch_req_0 : boolean;
  signal if_stmt_2679_branch_ack_1 : boolean;
  signal if_stmt_2679_branch_ack_0 : boolean;
  signal WPIPE_Block2_complete_2709_inst_req_0 : boolean;
  signal WPIPE_Block2_complete_2709_inst_ack_0 : boolean;
  signal WPIPE_Block2_complete_2709_inst_req_1 : boolean;
  signal WPIPE_Block2_complete_2709_inst_ack_1 : boolean;
  signal type_cast_2279_inst_req_0 : boolean;
  signal type_cast_2279_inst_ack_0 : boolean;
  signal type_cast_2279_inst_req_1 : boolean;
  signal type_cast_2279_inst_ack_1 : boolean;
  signal phi_stmt_2276_req_0 : boolean;
  signal phi_stmt_2282_req_0 : boolean;
  signal phi_stmt_2289_req_0 : boolean;
  signal type_cast_2281_inst_req_0 : boolean;
  signal type_cast_2281_inst_ack_0 : boolean;
  signal type_cast_2281_inst_req_1 : boolean;
  signal type_cast_2281_inst_ack_1 : boolean;
  signal phi_stmt_2276_req_1 : boolean;
  signal type_cast_2701_inst_ack_0 : boolean;
  signal type_cast_2701_inst_req_1 : boolean;
  signal type_cast_2701_inst_ack_1 : boolean;
  signal phi_stmt_2698_req_0 : boolean;
  signal phi_stmt_2686_ack_0 : boolean;
  signal phi_stmt_2692_ack_0 : boolean;
  signal phi_stmt_2698_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_C_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_C_CP_5741_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_C_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_C_CP_5741_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_C_CP_5741_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_C_CP_5741_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_C_CP_5741: Block -- control-path 
    signal zeropad3D_C_CP_5741_elements: BooleanArray(138 downto 0);
    -- 
  begin -- 
    zeropad3D_C_CP_5741_elements(0) <= zeropad3D_C_CP_5741_start;
    zeropad3D_C_CP_5741_symbol <= zeropad3D_C_CP_5741_elements(92);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2086/$entry
      -- CP-element group 0: 	 branch_block_stmt_2086/branch_block_stmt_2086__entry__
      -- CP-element group 0: 	 branch_block_stmt_2086/assign_stmt_2089__entry__
      -- CP-element group 0: 	 branch_block_stmt_2086/assign_stmt_2089/$entry
      -- CP-element group 0: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Sample/rr
      -- 
    rr_5819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(0), ack => RPIPE_Block2_starting_2088_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	138 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	100 
    -- CP-element group 1: 	102 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	105 
    -- CP-element group 1: 	106 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/merge_stmt_2685__exit__
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/$entry
      -- CP-element group 1: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/$entry
      -- 
    rr_7060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(1), ack => type_cast_2295_inst_req_0); -- 
    cr_7065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(1), ack => type_cast_2295_inst_req_1); -- 
    cr_7042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(1), ack => type_cast_2288_inst_req_1); -- 
    rr_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(1), ack => type_cast_2288_inst_req_0); -- 
    rr_7014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(1), ack => type_cast_2281_inst_req_0); -- 
    cr_7019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(1), ack => type_cast_2281_inst_req_1); -- 
    zeropad3D_C_CP_5741_elements(1) <= zeropad3D_C_CP_5741_elements(138);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Update/cr
      -- 
    ra_5820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_2088_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(2)); -- 
    cr_5824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(2), ack => RPIPE_Block2_starting_2088_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	17 
    -- CP-element group 3: 	19 
    -- CP-element group 3: 	13 
    -- CP-element group 3: 	10 
    -- CP-element group 3: 	16 
    -- CP-element group 3: 	14 
    -- CP-element group 3: 	15 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	7 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	9 
    -- CP-element group 3:  members (155) 
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2089__exit__
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273__entry__
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2089/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2089/RPIPE_Block2_starting_2088_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Update/cr
      -- 
    ca_5825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_2088_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(3)); -- 
    cr_5969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2126_load_0_req_1); -- 
    rr_6008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2138_load_0_req_0); -- 
    rr_5958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2126_load_0_req_0); -- 
    cr_6019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2138_load_0_req_1); -- 
    cr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => type_cast_2111_inst_req_1); -- 
    rr_6058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2150_load_0_req_0); -- 
    rr_5908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => LOAD_pad_2114_load_0_req_0); -- 
    rr_5861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2101_load_0_req_0); -- 
    cr_6069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2150_load_0_req_1); -- 
    cr_5919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => LOAD_pad_2114_load_0_req_1); -- 
    rr_6108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2162_load_0_req_0); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2101_load_0_req_1); -- 
    cr_6119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => ptr_deref_2162_load_0_req_1); -- 
    cr_6138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(3), ack => type_cast_2216_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/word_access_start/$exit
      -- CP-element group 4: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Sample/word_access_start/word_0/ra
      -- CP-element group 4: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_sample_completed_
      -- 
    ra_5862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2101_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (12) 
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/ptr_deref_2101_Merge/merge_ack
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/ptr_deref_2101_Merge/merge_req
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/ptr_deref_2101_Merge/$exit
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/ptr_deref_2101_Merge/$entry
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/word_access_complete/word_0/ca
      -- CP-element group 5: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2101_Update/$exit
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2101_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(5)); -- 
    rr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(5), ack => type_cast_2111_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_sample_completed_
      -- 
    ra_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2111_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	3 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2111_Update/ca
      -- 
    ca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2111_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Sample/word_access_start/$exit
      -- 
    ra_5909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2114_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	3 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	18 
    -- CP-element group 9:  members (12) 
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/LOAD_pad_2114_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/LOAD_pad_2114_Merge/merge_ack
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/LOAD_pad_2114_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/LOAD_pad_2114_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/LOAD_pad_2114_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Sample/rr
      -- 
    ca_5920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2114_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(9)); -- 
    rr_6133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(9), ack => type_cast_2216_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/word_access_start/$exit
      -- CP-element group 10: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Sample/word_access_start/word_0/ra
      -- 
    ra_5959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2126_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	20 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/word_access_complete/$exit
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/word_access_complete/word_0/ca
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/ptr_deref_2126_Merge/$entry
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/ptr_deref_2126_Merge/$exit
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/ptr_deref_2126_Merge/merge_req
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/ptr_deref_2126_Merge/merge_ack
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2126_Update/word_access_complete/word_0/$exit
      -- 
    ca_5970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2126_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/word_access_start/$exit
      -- CP-element group 12: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/word_access_start/word_0/ra
      -- CP-element group 12: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Sample/word_access_start/word_0/$exit
      -- 
    ra_6009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2138_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	20 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/ptr_deref_2138_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/ptr_deref_2138_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/ptr_deref_2138_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2138_Update/ptr_deref_2138_Merge/merge_ack
      -- 
    ca_6020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2138_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	3 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/word_access_start/word_0/ra
      -- CP-element group 14: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_sample_completed_
      -- 
    ra_6059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2150_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/ptr_deref_2150_Merge/merge_ack
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/ptr_deref_2150_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/ptr_deref_2150_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/ptr_deref_2150_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2150_Update/word_access_complete/word_0/ca
      -- 
    ca_6070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2150_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Sample/word_access_start/word_0/ra
      -- 
    ra_6109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2162_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/ptr_deref_2162_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/ptr_deref_2162_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/ptr_deref_2162_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/ptr_deref_2162_Update/ptr_deref_2162_Merge/merge_ack
      -- 
    ca_6120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2162_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	9 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Sample/ra
      -- 
    ra_6134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2216_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	3 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/type_cast_2216_Update/ca
      -- 
    ca_6139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2216_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  place  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	19 
    -- CP-element group 20: 	13 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	93 
    -- CP-element group 20: 	94 
    -- CP-element group 20: 	96 
    -- CP-element group 20: 	97 
    -- CP-element group 20:  members (16) 
      -- CP-element group 20: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273__exit__
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody
      -- CP-element group 20: 	 branch_block_stmt_2086/assign_stmt_2098_to_assign_stmt_2273/$exit
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2282/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2289/$entry
      -- CP-element group 20: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$entry
      -- 
    rr_6972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(20), ack => type_cast_2279_inst_req_0); -- 
    cr_6977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(20), ack => type_cast_2279_inst_req_1); -- 
    zeropad3D_C_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(11) & zeropad3D_C_CP_5741_elements(17) & zeropad3D_C_CP_5741_elements(19) & zeropad3D_C_CP_5741_elements(13) & zeropad3D_C_CP_5741_elements(15) & zeropad3D_C_CP_5741_elements(7);
      gj_zeropad3D_C_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	113 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Sample/ra
      -- 
    ra_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(21)); -- 
    -- CP-element group 22:  branch  transition  place  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	113 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (13) 
      -- CP-element group 22: 	 branch_block_stmt_2086/R_cmp_2310_place
      -- CP-element group 22: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308__exit__
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309__entry__
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309_dead_link/$entry
      -- CP-element group 22: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/$exit
      -- CP-element group 22: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309_eval_test/$entry
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309_eval_test/$exit
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309_eval_test/branch_req
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309_if_link/$entry
      -- CP-element group 22: 	 branch_block_stmt_2086/if_stmt_2309_else_link/$entry
      -- 
    ca_6156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(22)); -- 
    branch_req_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(22), ack => if_stmt_2309_branch_req_0); -- 
    -- CP-element group 23:  transition  place  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	114 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_2086/whilex_xbody_ifx_xthen
      -- CP-element group 23: 	 branch_block_stmt_2086/if_stmt_2309_if_link/$exit
      -- CP-element group 23: 	 branch_block_stmt_2086/if_stmt_2309_if_link/if_choice_transition
      -- CP-element group 23: 	 branch_block_stmt_2086/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_2086/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- 
    if_choice_transition_6169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2309_branch_ack_1, ack => zeropad3D_C_CP_5741_elements(23)); -- 
    -- CP-element group 24:  merge  transition  place  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (11) 
      -- CP-element group 24: 	 branch_block_stmt_2086/merge_stmt_2315_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_2086/merge_stmt_2315_PhiAck/dummy
      -- CP-element group 24: 	 branch_block_stmt_2086/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 24: 	 branch_block_stmt_2086/merge_stmt_2315_PhiAck/$exit
      -- CP-element group 24: 	 branch_block_stmt_2086/merge_stmt_2315__exit__
      -- CP-element group 24: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337__entry__
      -- CP-element group 24: 	 branch_block_stmt_2086/if_stmt_2309_else_link/$exit
      -- CP-element group 24: 	 branch_block_stmt_2086/if_stmt_2309_else_link/else_choice_transition
      -- CP-element group 24: 	 branch_block_stmt_2086/merge_stmt_2315_PhiAck/$entry
      -- CP-element group 24: 	 branch_block_stmt_2086/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 24: 	 branch_block_stmt_2086/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- 
    else_choice_transition_6173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2309_branch_ack_0, ack => zeropad3D_C_CP_5741_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (27) 
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_update_start_
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_address_calculated
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_word_address_calculated
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_root_address_calculated
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_address_resized
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_addr_resize/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_addr_resize/$exit
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_addr_resize/base_resize_req
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_addr_resize/base_resize_ack
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_plus_offset/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_plus_offset/$exit
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_plus_offset/sum_rename_req
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_base_plus_offset/sum_rename_ack
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_word_addrgen/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_word_addrgen/$exit
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_word_addrgen/root_register_req
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_word_addrgen/root_register_ack
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/word_access_start/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/word_access_start/word_0/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/word_access_start/word_0/rr
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/word_access_complete/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/word_access_complete/word_0/$entry
      -- CP-element group 25: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/word_access_complete/word_0/cr
      -- 
    cr_6222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(25), ack => ptr_deref_2326_load_0_req_1); -- 
    rr_6211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(25), ack => ptr_deref_2326_load_0_req_0); -- 
    zeropad3D_C_CP_5741_elements(25) <= zeropad3D_C_CP_5741_elements(24);
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/word_access_start/$exit
      -- CP-element group 26: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/word_access_start/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Sample/word_access_start/word_0/ra
      -- 
    ra_6212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2326_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(26)); -- 
    -- CP-element group 27:  branch  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (19) 
      -- CP-element group 27: 	 branch_block_stmt_2086/R_cmp48_2339_place
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337__exit__
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338__entry__
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/$exit
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/word_access_complete/$exit
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/word_access_complete/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/word_access_complete/word_0/ca
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/ptr_deref_2326_Merge/$entry
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/ptr_deref_2326_Merge/$exit
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/ptr_deref_2326_Merge/merge_req
      -- CP-element group 27: 	 branch_block_stmt_2086/assign_stmt_2323_to_assign_stmt_2337/ptr_deref_2326_Update/ptr_deref_2326_Merge/merge_ack
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338_dead_link/$entry
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338_eval_test/$entry
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338_eval_test/$exit
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338_eval_test/branch_req
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338_if_link/$entry
      -- CP-element group 27: 	 branch_block_stmt_2086/if_stmt_2338_else_link/$entry
      -- 
    ca_6223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2326_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(27)); -- 
    branch_req_6236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(27), ack => if_stmt_2338_branch_req_0); -- 
    -- CP-element group 28:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (18) 
      -- CP-element group 28: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse50
      -- CP-element group 28: 	 branch_block_stmt_2086/merge_stmt_2344_PhiAck/dummy
      -- CP-element group 28: 	 branch_block_stmt_2086/merge_stmt_2344_PhiAck/$exit
      -- CP-element group 28: 	 branch_block_stmt_2086/merge_stmt_2344_PhiAck/$entry
      -- CP-element group 28: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse50_PhiReq/$exit
      -- CP-element group 28: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse50_PhiReq/$entry
      -- CP-element group 28: 	 branch_block_stmt_2086/merge_stmt_2344_PhiReqMerge
      -- CP-element group 28: 	 branch_block_stmt_2086/merge_stmt_2344__exit__
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356__entry__
      -- CP-element group 28: 	 branch_block_stmt_2086/if_stmt_2338_if_link/$exit
      -- CP-element group 28: 	 branch_block_stmt_2086/if_stmt_2338_if_link/if_choice_transition
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/$entry
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Update/cr
      -- 
    if_choice_transition_6241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2338_branch_ack_1, ack => zeropad3D_C_CP_5741_elements(28)); -- 
    rr_6258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(28), ack => type_cast_2348_inst_req_0); -- 
    cr_6263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(28), ack => type_cast_2348_inst_req_1); -- 
    -- CP-element group 29:  transition  place  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	114 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 29: 	 branch_block_stmt_2086/if_stmt_2338_else_link/$exit
      -- CP-element group 29: 	 branch_block_stmt_2086/if_stmt_2338_else_link/else_choice_transition
      -- CP-element group 29: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- CP-element group 29: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- 
    else_choice_transition_6245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2338_branch_ack_0, ack => zeropad3D_C_CP_5741_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Sample/ra
      -- 
    ra_6259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2348_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(30)); -- 
    -- CP-element group 31:  branch  transition  place  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	28 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (13) 
      -- CP-element group 31: 	 branch_block_stmt_2086/R_cmp55_2358_place
      -- CP-element group 31: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356__exit__
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357__entry__
      -- CP-element group 31: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/$exit
      -- CP-element group 31: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2086/assign_stmt_2349_to_assign_stmt_2356/type_cast_2348_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357_dead_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357_eval_test/$entry
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357_eval_test/$exit
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357_eval_test/branch_req
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357_if_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_2086/if_stmt_2357_else_link/$entry
      -- 
    ca_6264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2348_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(31)); -- 
    branch_req_6272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(31), ack => if_stmt_2357_branch_req_0); -- 
    -- CP-element group 32:  transition  place  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	114 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse50_ifx_xthen
      -- CP-element group 32: 	 branch_block_stmt_2086/if_stmt_2357_if_link/$exit
      -- CP-element group 32: 	 branch_block_stmt_2086/if_stmt_2357_if_link/if_choice_transition
      -- CP-element group 32: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse50_ifx_xthen_PhiReq/$exit
      -- CP-element group 32: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse50_ifx_xthen_PhiReq/$entry
      -- 
    if_choice_transition_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2357_branch_ack_1, ack => zeropad3D_C_CP_5741_elements(32)); -- 
    -- CP-element group 33:  merge  transition  place  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (11) 
      -- CP-element group 33: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse50_lorx_xlhsx_xfalse57
      -- CP-element group 33: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse50_lorx_xlhsx_xfalse57_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse50_lorx_xlhsx_xfalse57_PhiReq/$exit
      -- CP-element group 33: 	 branch_block_stmt_2086/merge_stmt_2363_PhiAck/$entry
      -- CP-element group 33: 	 branch_block_stmt_2086/merge_stmt_2363_PhiReqMerge
      -- CP-element group 33: 	 branch_block_stmt_2086/merge_stmt_2363_PhiAck/$exit
      -- CP-element group 33: 	 branch_block_stmt_2086/merge_stmt_2363_PhiAck/dummy
      -- CP-element group 33: 	 branch_block_stmt_2086/merge_stmt_2363__exit__
      -- CP-element group 33: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391__entry__
      -- CP-element group 33: 	 branch_block_stmt_2086/if_stmt_2357_else_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_2086/if_stmt_2357_else_link/else_choice_transition
      -- 
    else_choice_transition_6281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2357_branch_ack_0, ack => zeropad3D_C_CP_5741_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (27) 
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_word_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_root_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_address_resized
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_addr_resize/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_addr_resize/$exit
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_addr_resize/base_resize_req
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_addr_resize/base_resize_ack
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_plus_offset/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_plus_offset/$exit
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_plus_offset/sum_rename_req
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_base_plus_offset/sum_rename_ack
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_word_addrgen/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_word_addrgen/$exit
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_word_addrgen/root_register_req
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_word_addrgen/root_register_ack
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/word_access_start/word_0/rr
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/word_access_complete/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/word_access_complete/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/word_access_complete/word_0/cr
      -- 
    cr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(34), ack => ptr_deref_2374_load_0_req_1); -- 
    rr_6319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(34), ack => ptr_deref_2374_load_0_req_0); -- 
    zeropad3D_C_CP_5741_elements(34) <= zeropad3D_C_CP_5741_elements(33);
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/word_access_start/$exit
      -- CP-element group 35: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Sample/word_access_start/word_0/ra
      -- 
    ra_6320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2374_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (19) 
      -- CP-element group 36: 	 branch_block_stmt_2086/R_cmp65_2393_place
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391__exit__
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392__entry__
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/$exit
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/word_access_complete/word_0/ca
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/ptr_deref_2374_Merge/$entry
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/ptr_deref_2374_Merge/$exit
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/ptr_deref_2374_Merge/merge_req
      -- CP-element group 36: 	 branch_block_stmt_2086/assign_stmt_2371_to_assign_stmt_2391/ptr_deref_2374_Update/ptr_deref_2374_Merge/merge_ack
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2086/if_stmt_2392_else_link/$entry
      -- 
    ca_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2374_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(36)); -- 
    branch_req_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(36), ack => if_stmt_2392_branch_req_0); -- 
    -- CP-element group 37:  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	64 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	56 
    -- CP-element group 37: 	68 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	53 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	60 
    -- CP-element group 37: 	71 
    -- CP-element group 37:  members (46) 
      -- CP-element group 37: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse57_ifx_xelse
      -- CP-element group 37: 	 branch_block_stmt_2086/merge_stmt_2456_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_2086/merge_stmt_2456__exit__
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561__entry__
      -- CP-element group 37: 	 branch_block_stmt_2086/if_stmt_2392_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_2086/if_stmt_2392_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_2086/merge_stmt_2456_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_2086/merge_stmt_2456_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_2086/merge_stmt_2456_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse57_ifx_xelse_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse57_ifx_xelse_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_update_start
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Update/req
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_complete/req
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_update_start
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Update/req
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_complete/req
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/word_access_complete/word_0/cr
      -- 
    if_choice_transition_6349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2392_branch_ack_1, ack => zeropad3D_C_CP_5741_elements(37)); -- 
    rr_6507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => type_cast_2460_inst_req_0); -- 
    cr_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => type_cast_2460_inst_req_1); -- 
    cr_6526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => type_cast_2524_inst_req_1); -- 
    req_6557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => array_obj_ref_2530_index_offset_req_1); -- 
    req_6572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => addr_of_2531_final_reg_req_1); -- 
    cr_6617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => ptr_deref_2535_load_0_req_1); -- 
    cr_6636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => type_cast_2549_inst_req_1); -- 
    req_6667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => array_obj_ref_2555_index_offset_req_1); -- 
    req_6682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => addr_of_2556_final_reg_req_1); -- 
    cr_6732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(37), ack => ptr_deref_2559_store_0_req_1); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	114 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse57_ifx_xthen
      -- CP-element group 38: 	 branch_block_stmt_2086/if_stmt_2392_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_2086/if_stmt_2392_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse57_ifx_xthen_PhiReq/$exit
      -- CP-element group 38: 	 branch_block_stmt_2086/lorx_xlhsx_xfalse57_ifx_xthen_PhiReq/$entry
      -- 
    else_choice_transition_6353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2392_branch_ack_0, ack => zeropad3D_C_CP_5741_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	114 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Sample/ra
      -- 
    ra_6367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2402_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	114 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Update/ca
      -- 
    ca_6372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2402_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	114 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Sample/ra
      -- 
    ra_6381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2407_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	114 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Update/ca
      -- 
    ca_6386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2407_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: 	40 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Sample/rr
      -- 
    rr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(43), ack => type_cast_2441_inst_req_0); -- 
    zeropad3D_C_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(42) & zeropad3D_C_CP_5741_elements(40);
      gj_zeropad3D_C_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Sample/ra
      -- 
    ra_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	114 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Sample/req
      -- 
    ca_6400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(45)); -- 
    req_6425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(45), ack => array_obj_ref_2447_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	52 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Sample/ack
      -- 
    ack_6426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2447_index_offset_ack_0, ack => zeropad3D_C_CP_5741_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	114 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_request/req
      -- 
    ack_6431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2447_index_offset_ack_1, ack => zeropad3D_C_CP_5741_elements(47)); -- 
    req_6440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(47), ack => addr_of_2448_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_request/ack
      -- 
    ack_6441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2448_final_reg_ack_0, ack => zeropad3D_C_CP_5741_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	114 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (28) 
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/ptr_deref_2451_Split/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/ptr_deref_2451_Split/$exit
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/ptr_deref_2451_Split/split_req
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/ptr_deref_2451_Split/split_ack
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/word_access_start/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/word_access_start/word_0/$entry
      -- CP-element group 49: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/word_access_start/word_0/rr
      -- 
    ack_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2448_final_reg_ack_1, ack => zeropad3D_C_CP_5741_elements(49)); -- 
    rr_6484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(49), ack => ptr_deref_2451_store_0_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Sample/word_access_start/word_0/ra
      -- 
    ra_6485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2451_store_0_ack_0, ack => zeropad3D_C_CP_5741_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	114 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/word_access_complete/word_0/ca
      -- 
    ca_6496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2451_store_0_ack_1, ack => zeropad3D_C_CP_5741_elements(51)); -- 
    -- CP-element group 52:  join  transition  place  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	46 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	115 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454__exit__
      -- CP-element group 52: 	 branch_block_stmt_2086/ifx_xthen_ifx_xend
      -- CP-element group 52: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/$exit
      -- CP-element group 52: 	 branch_block_stmt_2086/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_2086/ifx_xthen_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_C_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(46) & zeropad3D_C_CP_5741_elements(51);
      gj_zeropad3D_C_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	37 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Sample/ra
      -- 
    ra_6508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	63 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2460_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Sample/rr
      -- 
    ca_6513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(54)); -- 
    rr_6631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(54), ack => type_cast_2549_inst_req_0); -- 
    rr_6521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(54), ack => type_cast_2524_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Sample/ra
      -- 
    ra_6522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2524_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	37 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (16) 
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2524_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Sample/req
      -- 
    ca_6527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2524_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(56)); -- 
    req_6552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(56), ack => array_obj_ref_2530_index_offset_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	72 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Sample/ack
      -- 
    ack_6553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2530_index_offset_ack_0, ack => zeropad3D_C_CP_5741_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2530_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_request/req
      -- 
    ack_6558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2530_index_offset_ack_1, ack => zeropad3D_C_CP_5741_elements(58)); -- 
    req_6567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(58), ack => addr_of_2531_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_request/ack
      -- 
    ack_6568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2531_final_reg_ack_0, ack => zeropad3D_C_CP_5741_elements(59)); -- 
    -- CP-element group 60:  join  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	37 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2531_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_word_addrgen/root_register_ack
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/word_access_start/$entry
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/word_access_start/word_0/$entry
      -- CP-element group 60: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/word_access_start/word_0/rr
      -- 
    ack_6573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2531_final_reg_ack_1, ack => zeropad3D_C_CP_5741_elements(60)); -- 
    rr_6606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(60), ack => ptr_deref_2535_load_0_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/word_access_start/$exit
      -- CP-element group 61: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/word_access_start/word_0/$exit
      -- CP-element group 61: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Sample/word_access_start/word_0/ra
      -- 
    ra_6607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2535_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	69 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/word_access_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/word_access_complete/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/word_access_complete/word_0/ca
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/ptr_deref_2535_Merge/$entry
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/ptr_deref_2535_Merge/$exit
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/ptr_deref_2535_Merge/merge_req
      -- CP-element group 62: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2535_Update/ptr_deref_2535_Merge/merge_ack
      -- 
    ca_6618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2535_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	54 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Sample/ra
      -- 
    ra_6632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	37 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (16) 
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/type_cast_2549_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_resized_1
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_scaled_1
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_computed_1
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_resize_1/$entry
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_resize_1/$exit
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_resize_1/index_resize_req
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_resize_1/index_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_scale_1/$entry
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_scale_1/$exit
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_scale_1/scale_rename_req
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_index_scale_1/scale_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Sample/req
      -- 
    ca_6637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(64)); -- 
    req_6662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(64), ack => array_obj_ref_2555_index_offset_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	72 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_sample_complete
      -- CP-element group 65: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Sample/ack
      -- 
    ack_6663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2555_index_offset_ack_0, ack => zeropad3D_C_CP_5741_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (11) 
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_root_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_offset_calculated
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_final_index_sum_regn_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_base_plus_offset/$entry
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_base_plus_offset/$exit
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_base_plus_offset/sum_rename_req
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/array_obj_ref_2555_base_plus_offset/sum_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_request/$entry
      -- CP-element group 66: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_request/req
      -- 
    ack_6668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2555_index_offset_ack_1, ack => zeropad3D_C_CP_5741_elements(66)); -- 
    req_6677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(66), ack => addr_of_2556_final_reg_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_request/$exit
      -- CP-element group 67: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_request/ack
      -- 
    ack_6678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2556_final_reg_ack_0, ack => zeropad3D_C_CP_5741_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	37 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (19) 
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_complete/$exit
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/addr_of_2556_complete/ack
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_word_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_address_resized
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_addr_resize/$entry
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_addr_resize/$exit
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_addr_resize/base_resize_req
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_addr_resize/base_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_word_addrgen/$entry
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_word_addrgen/$exit
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_word_addrgen/root_register_req
      -- CP-element group 68: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_word_addrgen/root_register_ack
      -- 
    ack_6683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2556_final_reg_ack_1, ack => zeropad3D_C_CP_5741_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: 	62 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (9) 
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/ptr_deref_2559_Split/$entry
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/ptr_deref_2559_Split/$exit
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/ptr_deref_2559_Split/split_req
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/ptr_deref_2559_Split/split_ack
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/word_access_start/$entry
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/word_access_start/word_0/$entry
      -- CP-element group 69: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/word_access_start/word_0/rr
      -- 
    rr_6721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(69), ack => ptr_deref_2559_store_0_req_0); -- 
    zeropad3D_C_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(68) & zeropad3D_C_CP_5741_elements(62);
      gj_zeropad3D_C_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/word_access_start/$exit
      -- CP-element group 70: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/word_access_start/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Sample/word_access_start/word_0/ra
      -- 
    ra_6722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2559_store_0_ack_0, ack => zeropad3D_C_CP_5741_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	37 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/word_access_complete/$exit
      -- CP-element group 71: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/word_access_complete/word_0/$exit
      -- CP-element group 71: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/ptr_deref_2559_Update/word_access_complete/word_0/ca
      -- 
    ca_6733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2559_store_0_ack_1, ack => zeropad3D_C_CP_5741_elements(71)); -- 
    -- CP-element group 72:  join  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	65 
    -- CP-element group 72: 	57 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	115 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561__exit__
      -- CP-element group 72: 	 branch_block_stmt_2086/ifx_xelse_ifx_xend
      -- CP-element group 72: 	 branch_block_stmt_2086/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_2086/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2086/assign_stmt_2461_to_assign_stmt_2561/$exit
      -- 
    zeropad3D_C_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(65) & zeropad3D_C_CP_5741_elements(57) & zeropad3D_C_CP_5741_elements(71);
      gj_zeropad3D_C_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	115 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Sample/ra
      -- 
    ra_6745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2567_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	115 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581__exit__
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582__entry__
      -- CP-element group 74: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/$exit
      -- CP-element group 74: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2086/R_cmp134_2583_place
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2086/if_stmt_2582_else_link/$entry
      -- 
    ca_6750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2567_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(74)); -- 
    branch_req_6758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(74), ack => if_stmt_2582_branch_req_0); -- 
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	124 
    -- CP-element group 75: 	125 
    -- CP-element group 75: 	127 
    -- CP-element group 75: 	128 
    -- CP-element group 75: 	130 
    -- CP-element group 75: 	131 
    -- CP-element group 75:  members (40) 
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/merge_stmt_2588_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2086/merge_stmt_2588__exit__
      -- CP-element group 75: 	 branch_block_stmt_2086/assign_stmt_2594__entry__
      -- CP-element group 75: 	 branch_block_stmt_2086/assign_stmt_2594__exit__
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/merge_stmt_2588_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_2086/merge_stmt_2588_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2086/merge_stmt_2588_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xend_ifx_xthen136_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xend_ifx_xthen136_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/if_stmt_2582_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2086/if_stmt_2582_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xend_ifx_xthen136
      -- CP-element group 75: 	 branch_block_stmt_2086/assign_stmt_2594/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/assign_stmt_2594/$exit
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2582_branch_ack_1, ack => zeropad3D_C_CP_5741_elements(75)); -- 
    rr_7296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(75), ack => type_cast_2701_inst_req_0); -- 
    rr_7250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(75), ack => type_cast_2689_inst_req_0); -- 
    cr_7278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(75), ack => type_cast_2695_inst_req_1); -- 
    cr_7255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(75), ack => type_cast_2689_inst_req_1); -- 
    rr_7273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(75), ack => type_cast_2695_inst_req_0); -- 
    cr_7301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(75), ack => type_cast_2701_inst_req_1); -- 
    -- CP-element group 76:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76: 	79 
    -- CP-element group 76: 	80 
    -- CP-element group 76: 	83 
    -- CP-element group 76: 	85 
    -- CP-element group 76: 	86 
    -- CP-element group 76: 	87 
    -- CP-element group 76:  members (76) 
      -- CP-element group 76: 	 branch_block_stmt_2086/merge_stmt_2596_PhiAck/dummy
      -- CP-element group 76: 	 branch_block_stmt_2086/merge_stmt_2596_PhiAck/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/merge_stmt_2596_PhiAck/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/merge_stmt_2596_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_2086/merge_stmt_2596__exit__
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678__entry__
      -- CP-element group 76: 	 branch_block_stmt_2086/ifx_xend_ifx_xelse141_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/ifx_xend_ifx_xelse141_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/if_stmt_2582_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/if_stmt_2582_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2086/ifx_xend_ifx_xelse141
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_update_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_update_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_word_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_root_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_address_resized
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_addr_resize/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_addr_resize/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_addr_resize/base_resize_req
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_addr_resize/base_resize_ack
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_plus_offset/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_plus_offset/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_plus_offset/sum_rename_req
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_base_plus_offset/sum_rename_ack
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_word_addrgen/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_word_addrgen/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_word_addrgen/root_register_req
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_word_addrgen/root_register_ack
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/word_access_start/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/word_access_start/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/word_access_start/word_0/rr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/word_access_complete/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/word_access_complete/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/word_access_complete/word_0/cr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_update_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_update_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_update_start_
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_word_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_root_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_address_resized
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_addr_resize/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_addr_resize/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_addr_resize/base_resize_req
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_addr_resize/base_resize_ack
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_plus_offset/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_plus_offset/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_plus_offset/sum_rename_req
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_base_plus_offset/sum_rename_ack
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_word_addrgen/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_word_addrgen/$exit
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_word_addrgen/root_register_req
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_word_addrgen/root_register_ack
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/word_access_start/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/word_access_start/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/word_access_start/word_0/rr
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/word_access_complete/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/word_access_complete/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2582_branch_ack_0, ack => zeropad3D_C_CP_5741_elements(76)); -- 
    rr_6783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => type_cast_2606_inst_req_0); -- 
    cr_6788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => type_cast_2606_inst_req_1); -- 
    rr_6822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => ptr_deref_2618_load_0_req_0); -- 
    cr_6833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => ptr_deref_2618_load_0_req_1); -- 
    cr_6852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => type_cast_2638_inst_req_1); -- 
    cr_6866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => type_cast_2655_inst_req_1); -- 
    rr_6900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => ptr_deref_2667_load_0_req_0); -- 
    cr_6911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(76), ack => ptr_deref_2667_load_0_req_1); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Sample/ra
      -- 
    ra_6784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2606_Update/ca
      -- 
    ca_6789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	76 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/word_access_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/word_access_start/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Sample/word_access_start/word_0/ra
      -- 
    ra_6823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2618_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	76 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/word_access_complete/word_0/ca
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/ptr_deref_2618_Merge/$entry
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/ptr_deref_2618_Merge/$exit
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/ptr_deref_2618_Merge/merge_req
      -- CP-element group 80: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2618_Update/ptr_deref_2618_Merge/merge_ack
      -- 
    ca_6834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2618_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Sample/rr
      -- 
    rr_6847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(81), ack => type_cast_2638_inst_req_0); -- 
    zeropad3D_C_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(78) & zeropad3D_C_CP_5741_elements(80);
      gj_zeropad3D_C_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Sample/ra
      -- 
    ra_6848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2638_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	76 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2638_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Sample/rr
      -- 
    ca_6853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2638_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(83)); -- 
    rr_6861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(83), ack => type_cast_2655_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Sample/ra
      -- 
    ra_6862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	76 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	88 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/type_cast_2655_Update/ca
      -- 
    ca_6867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	76 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/word_access_start/$exit
      -- CP-element group 86: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/word_access_start/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Sample/word_access_start/word_0/ra
      -- 
    ra_6901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_load_0_ack_0, ack => zeropad3D_C_CP_5741_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	76 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/word_access_complete/$exit
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/word_access_complete/word_0/$exit
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/word_access_complete/word_0/ca
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/ptr_deref_2667_Merge/$entry
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/ptr_deref_2667_Merge/$exit
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/ptr_deref_2667_Merge/merge_req
      -- CP-element group 87: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/ptr_deref_2667_Update/ptr_deref_2667_Merge/merge_ack
      -- 
    ca_6912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2667_load_0_ack_1, ack => zeropad3D_C_CP_5741_elements(87)); -- 
    -- CP-element group 88:  branch  join  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	85 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (10) 
      -- CP-element group 88: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678__exit__
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679__entry__
      -- CP-element group 88: 	 branch_block_stmt_2086/assign_stmt_2602_to_assign_stmt_2678/$exit
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679_dead_link/$entry
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679_eval_test/$entry
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679_eval_test/$exit
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679_eval_test/branch_req
      -- CP-element group 88: 	 branch_block_stmt_2086/R_cmp164_2680_place
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679_if_link/$entry
      -- CP-element group 88: 	 branch_block_stmt_2086/if_stmt_2679_else_link/$entry
      -- 
    branch_req_6925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(88), ack => if_stmt_2679_branch_req_0); -- 
    zeropad3D_C_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(85) & zeropad3D_C_CP_5741_elements(87);
      gj_zeropad3D_C_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (15) 
      -- CP-element group 89: 	 branch_block_stmt_2086/merge_stmt_2707__exit__
      -- CP-element group 89: 	 branch_block_stmt_2086/assign_stmt_2711__entry__
      -- CP-element group 89: 	 branch_block_stmt_2086/if_stmt_2679_if_link/$exit
      -- CP-element group 89: 	 branch_block_stmt_2086/if_stmt_2679_if_link/if_choice_transition
      -- CP-element group 89: 	 branch_block_stmt_2086/ifx_xelse141_whilex_xend
      -- CP-element group 89: 	 branch_block_stmt_2086/assign_stmt_2711/$entry
      -- CP-element group 89: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Sample/req
      -- CP-element group 89: 	 branch_block_stmt_2086/ifx_xelse141_whilex_xend_PhiReq/$entry
      -- CP-element group 89: 	 branch_block_stmt_2086/ifx_xelse141_whilex_xend_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2086/merge_stmt_2707_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2086/merge_stmt_2707_PhiAck/$entry
      -- CP-element group 89: 	 branch_block_stmt_2086/merge_stmt_2707_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_2086/merge_stmt_2707_PhiAck/dummy
      -- 
    if_choice_transition_6930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2679_branch_ack_1, ack => zeropad3D_C_CP_5741_elements(89)); -- 
    req_6947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(89), ack => WPIPE_Block2_complete_2709_inst_req_0); -- 
    -- CP-element group 90:  fork  transition  place  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	116 
    -- CP-element group 90: 	117 
    -- CP-element group 90: 	119 
    -- CP-element group 90: 	120 
    -- CP-element group 90: 	122 
    -- CP-element group 90:  members (22) 
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Update/cr
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2698/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Update/cr
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/$entry
      -- CP-element group 90: 	 branch_block_stmt_2086/if_stmt_2679_else_link/$exit
      -- CP-element group 90: 	 branch_block_stmt_2086/if_stmt_2679_else_link/else_choice_transition
      -- CP-element group 90: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172
      -- 
    else_choice_transition_6934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2679_branch_ack_0, ack => zeropad3D_C_CP_5741_elements(90)); -- 
    cr_7221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(90), ack => type_cast_2697_inst_req_1); -- 
    rr_7216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(90), ack => type_cast_2697_inst_req_0); -- 
    cr_7198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(90), ack => type_cast_2691_inst_req_1); -- 
    rr_7193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(90), ack => type_cast_2691_inst_req_0); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Update/req
      -- 
    ack_6948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_complete_2709_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(91)); -- 
    req_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(91), ack => WPIPE_Block2_complete_2709_inst_req_1); -- 
    -- CP-element group 92:  transition  place  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (16) 
      -- CP-element group 92: 	 $exit
      -- CP-element group 92: 	 branch_block_stmt_2086/$exit
      -- CP-element group 92: 	 branch_block_stmt_2086/branch_block_stmt_2086__exit__
      -- CP-element group 92: 	 branch_block_stmt_2086/assign_stmt_2711__exit__
      -- CP-element group 92: 	 branch_block_stmt_2086/return__
      -- CP-element group 92: 	 branch_block_stmt_2086/merge_stmt_2713__exit__
      -- CP-element group 92: 	 branch_block_stmt_2086/assign_stmt_2711/$exit
      -- CP-element group 92: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2086/assign_stmt_2711/WPIPE_Block2_complete_2709_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_2086/return___PhiReq/$entry
      -- CP-element group 92: 	 branch_block_stmt_2086/return___PhiReq/$exit
      -- CP-element group 92: 	 branch_block_stmt_2086/merge_stmt_2713_PhiReqMerge
      -- CP-element group 92: 	 branch_block_stmt_2086/merge_stmt_2713_PhiAck/$entry
      -- CP-element group 92: 	 branch_block_stmt_2086/merge_stmt_2713_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_2086/merge_stmt_2713_PhiAck/dummy
      -- 
    ack_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_complete_2709_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	20 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/ra
      -- 
    ra_6973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	20 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/ca
      -- 
    ca_6978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/$exit
      -- CP-element group 95: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/$exit
      -- CP-element group 95: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_req
      -- 
    phi_stmt_2276_req_6979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2276_req_6979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(95), ack => phi_stmt_2276_req_0); -- 
    zeropad3D_C_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(93) & zeropad3D_C_CP_5741_elements(94);
      gj_zeropad3D_C_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  output  delay-element  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	20 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2282/$exit
      -- CP-element group 96: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2286_konst_delay_trans
      -- CP-element group 96: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_req
      -- 
    phi_stmt_2282_req_6987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2282_req_6987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(96), ack => phi_stmt_2282_req_0); -- 
    -- Element group zeropad3D_C_CP_5741_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_5741_elements(20), ack => zeropad3D_C_CP_5741_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  transition  output  delay-element  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	20 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2289/$exit
      -- CP-element group 97: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2293_konst_delay_trans
      -- CP-element group 97: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_req
      -- 
    phi_stmt_2289_req_6995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2289_req_6995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(97), ack => phi_stmt_2289_req_0); -- 
    -- Element group zeropad3D_C_CP_5741_elements(97) is a control-delay.
    cp_element_97_delay: control_delay_element  generic map(name => " 97_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_5741_elements(20), ack => zeropad3D_C_CP_5741_elements(97), clk => clk, reset =>reset);
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: 	96 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	109 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2086/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(95) & zeropad3D_C_CP_5741_elements(96) & zeropad3D_C_CP_5741_elements(97);
      gj_zeropad3D_C_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/ra
      -- 
    ra_7015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2281_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/ca
      -- 
    ca_7020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2281_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/$exit
      -- CP-element group 101: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/$exit
      -- CP-element group 101: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2276/phi_stmt_2276_req
      -- 
    phi_stmt_2276_req_7021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2276_req_7021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(101), ack => phi_stmt_2276_req_1); -- 
    zeropad3D_C_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(99) & zeropad3D_C_CP_5741_elements(100);
      gj_zeropad3D_C_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/$exit
      -- 
    ra_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/ca
      -- CP-element group 103: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/$exit
      -- 
    ca_7043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_req
      -- CP-element group 104: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/$exit
      -- CP-element group 104: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/$exit
      -- CP-element group 104: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/$exit
      -- 
    phi_stmt_2282_req_7044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2282_req_7044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(104), ack => phi_stmt_2282_req_1); -- 
    zeropad3D_C_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(102) & zeropad3D_C_CP_5741_elements(103);
      gj_zeropad3D_C_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	1 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/$exit
      -- 
    ra_7061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/ca
      -- 
    ca_7066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/$exit
      -- CP-element group 107: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/$exit
      -- CP-element group 107: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_req
      -- 
    phi_stmt_2289_req_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2289_req_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(107), ack => phi_stmt_2289_req_1); -- 
    zeropad3D_C_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(105) & zeropad3D_C_CP_5741_elements(106);
      gj_zeropad3D_C_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2086/ifx_xend172_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(101) & zeropad3D_C_CP_5741_elements(104) & zeropad3D_C_CP_5741_elements(107);
      gj_zeropad3D_C_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	98 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2086/merge_stmt_2275_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_2086/merge_stmt_2275_PhiAck/$entry
      -- 
    zeropad3D_C_CP_5741_elements(109) <= OrReduce(zeropad3D_C_CP_5741_elements(98) & zeropad3D_C_CP_5741_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_2086/merge_stmt_2275_PhiAck/phi_stmt_2276_ack
      -- 
    phi_stmt_2276_ack_7072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2276_ack_0, ack => zeropad3D_C_CP_5741_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2086/merge_stmt_2275_PhiAck/phi_stmt_2282_ack
      -- 
    phi_stmt_2282_ack_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2282_ack_0, ack => zeropad3D_C_CP_5741_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2086/merge_stmt_2275_PhiAck/phi_stmt_2289_ack
      -- 
    phi_stmt_2289_ack_7074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2289_ack_0, ack => zeropad3D_C_CP_5741_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	21 
    -- CP-element group 113: 	22 
    -- CP-element group 113:  members (10) 
      -- CP-element group 113: 	 branch_block_stmt_2086/merge_stmt_2275__exit__
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308__entry__
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/$entry
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_update_start_
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_2086/assign_stmt_2301_to_assign_stmt_2308/type_cast_2300_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_2086/merge_stmt_2275_PhiAck/$exit
      -- 
    rr_6150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(113), ack => type_cast_2300_inst_req_0); -- 
    cr_6155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(113), ack => type_cast_2300_inst_req_1); -- 
    zeropad3D_C_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(110) & zeropad3D_C_CP_5741_elements(111) & zeropad3D_C_CP_5741_elements(112);
      gj_zeropad3D_C_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  merge  fork  transition  place  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	38 
    -- CP-element group 114: 	29 
    -- CP-element group 114: 	32 
    -- CP-element group 114: 	23 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	49 
    -- CP-element group 114: 	42 
    -- CP-element group 114: 	41 
    -- CP-element group 114: 	39 
    -- CP-element group 114: 	40 
    -- CP-element group 114: 	47 
    -- CP-element group 114: 	45 
    -- CP-element group 114: 	51 
    -- CP-element group 114:  members (33) 
      -- CP-element group 114: 	 branch_block_stmt_2086/merge_stmt_2398_PhiReqMerge
      -- CP-element group 114: 	 branch_block_stmt_2086/merge_stmt_2398__exit__
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454__entry__
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2402_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2407_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/type_cast_2441_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_update_start
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/array_obj_ref_2447_final_index_sum_regn_Update/req
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/addr_of_2448_complete/req
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/word_access_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/word_access_complete/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_2086/assign_stmt_2403_to_assign_stmt_2454/ptr_deref_2451_Update/word_access_complete/word_0/cr
      -- CP-element group 114: 	 branch_block_stmt_2086/merge_stmt_2398_PhiAck/dummy
      -- CP-element group 114: 	 branch_block_stmt_2086/merge_stmt_2398_PhiAck/$exit
      -- CP-element group 114: 	 branch_block_stmt_2086/merge_stmt_2398_PhiAck/$entry
      -- 
    rr_6366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => type_cast_2402_inst_req_0); -- 
    cr_6371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => type_cast_2402_inst_req_1); -- 
    rr_6380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => type_cast_2407_inst_req_0); -- 
    cr_6385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => type_cast_2407_inst_req_1); -- 
    cr_6399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => type_cast_2441_inst_req_1); -- 
    req_6430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => array_obj_ref_2447_index_offset_req_1); -- 
    req_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => addr_of_2448_final_reg_req_1); -- 
    cr_6495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(114), ack => ptr_deref_2451_store_0_req_1); -- 
    zeropad3D_C_CP_5741_elements(114) <= OrReduce(zeropad3D_C_CP_5741_elements(38) & zeropad3D_C_CP_5741_elements(29) & zeropad3D_C_CP_5741_elements(32) & zeropad3D_C_CP_5741_elements(23));
    -- CP-element group 115:  merge  fork  transition  place  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	52 
    -- CP-element group 115: 	72 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	73 
    -- CP-element group 115: 	74 
    -- CP-element group 115:  members (13) 
      -- CP-element group 115: 	 branch_block_stmt_2086/merge_stmt_2563_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_2086/merge_stmt_2563__exit__
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581__entry__
      -- CP-element group 115: 	 branch_block_stmt_2086/merge_stmt_2563_PhiAck/dummy
      -- CP-element group 115: 	 branch_block_stmt_2086/merge_stmt_2563_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_2086/merge_stmt_2563_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/$entry
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_update_start_
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_2086/assign_stmt_2568_to_assign_stmt_2581/type_cast_2567_Update/cr
      -- 
    rr_6744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(115), ack => type_cast_2567_inst_req_0); -- 
    cr_6749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(115), ack => type_cast_2567_inst_req_1); -- 
    zeropad3D_C_CP_5741_elements(115) <= OrReduce(zeropad3D_C_CP_5741_elements(52) & zeropad3D_C_CP_5741_elements(72));
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	90 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Sample/$exit
      -- 
    ra_7194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2691_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	90 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/Update/$exit
      -- 
    ca_7199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2691_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/$exit
      -- CP-element group 118: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_req
      -- CP-element group 118: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2691/$exit
      -- 
    phi_stmt_2686_req_7200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2686_req_7200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(118), ack => phi_stmt_2686_req_1); -- 
    zeropad3D_C_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(116) & zeropad3D_C_CP_5741_elements(117);
      gj_zeropad3D_C_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	90 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Sample/$exit
      -- 
    ra_7217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	90 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/Update/ca
      -- 
    ca_7222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_req
      -- CP-element group 121: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2697/$exit
      -- CP-element group 121: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2692/$exit
      -- 
    phi_stmt_2692_req_7223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2692_req_7223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(121), ack => phi_stmt_2692_req_1); -- 
    zeropad3D_C_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(119) & zeropad3D_C_CP_5741_elements(120);
      gj_zeropad3D_C_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  output  delay-element  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	90 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2698/$exit
      -- CP-element group 122: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2704_konst_delay_trans
      -- CP-element group 122: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_req
      -- 
    phi_stmt_2698_req_7231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2698_req_7231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(122), ack => phi_stmt_2698_req_1); -- 
    -- Element group zeropad3D_C_CP_5741_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_5741_elements(90), ack => zeropad3D_C_CP_5741_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	134 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2086/ifx_xelse141_ifx_xend172_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(118) & zeropad3D_C_CP_5741_elements(121) & zeropad3D_C_CP_5741_elements(122);
      gj_zeropad3D_C_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	75 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Sample/ra
      -- 
    ra_7251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2689_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	75 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Update/ca
      -- CP-element group 125: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/Update/$exit
      -- 
    ca_7256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2689_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	133 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/$exit
      -- CP-element group 126: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/$exit
      -- CP-element group 126: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_req
      -- CP-element group 126: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2686/phi_stmt_2686_sources/type_cast_2689/SplitProtocol/$exit
      -- 
    phi_stmt_2686_req_7257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2686_req_7257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(126), ack => phi_stmt_2686_req_0); -- 
    zeropad3D_C_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(124) & zeropad3D_C_CP_5741_elements(125);
      gj_zeropad3D_C_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	75 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Sample/ra
      -- CP-element group 127: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Sample/$exit
      -- 
    ra_7274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	75 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Update/ca
      -- CP-element group 128: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/Update/$exit
      -- 
    ca_7279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_req
      -- CP-element group 129: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/$exit
      -- CP-element group 129: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/$exit
      -- CP-element group 129: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2692/phi_stmt_2692_sources/type_cast_2695/$exit
      -- 
    phi_stmt_2692_req_7280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2692_req_7280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(129), ack => phi_stmt_2692_req_0); -- 
    zeropad3D_C_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(127) & zeropad3D_C_CP_5741_elements(128);
      gj_zeropad3D_C_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	75 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Sample/ra
      -- 
    ra_7297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2701_inst_ack_0, ack => zeropad3D_C_CP_5741_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	75 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/Update/ca
      -- 
    ca_7302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2701_inst_ack_1, ack => zeropad3D_C_CP_5741_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/SplitProtocol/$exit
      -- CP-element group 132: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/$exit
      -- CP-element group 132: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/type_cast_2701/$exit
      -- CP-element group 132: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_sources/$exit
      -- CP-element group 132: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/phi_stmt_2698/phi_stmt_2698_req
      -- 
    phi_stmt_2698_req_7303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2698_req_7303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_5741_elements(132), ack => phi_stmt_2698_req_0); -- 
    zeropad3D_C_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(130) & zeropad3D_C_CP_5741_elements(131);
      gj_zeropad3D_C_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	126 
    -- CP-element group 133: 	129 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_2086/ifx_xthen136_ifx_xend172_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(126) & zeropad3D_C_CP_5741_elements(129) & zeropad3D_C_CP_5741_elements(132);
      gj_zeropad3D_C_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  merge  fork  transition  place  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	123 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2086/merge_stmt_2685_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_2086/merge_stmt_2685_PhiAck/$entry
      -- 
    zeropad3D_C_CP_5741_elements(134) <= OrReduce(zeropad3D_C_CP_5741_elements(123) & zeropad3D_C_CP_5741_elements(133));
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_2086/merge_stmt_2685_PhiAck/phi_stmt_2686_ack
      -- 
    phi_stmt_2686_ack_7308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2686_ack_0, ack => zeropad3D_C_CP_5741_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_2086/merge_stmt_2685_PhiAck/phi_stmt_2692_ack
      -- 
    phi_stmt_2692_ack_7309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2692_ack_0, ack => zeropad3D_C_CP_5741_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_2086/merge_stmt_2685_PhiAck/phi_stmt_2698_ack
      -- 
    phi_stmt_2698_ack_7310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2698_ack_0, ack => zeropad3D_C_CP_5741_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	1 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_2086/merge_stmt_2685_PhiAck/$exit
      -- 
    zeropad3D_C_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_5741_elements(135) & zeropad3D_C_CP_5741_elements(136) & zeropad3D_C_CP_5741_elements(137);
      gj_zeropad3D_C_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_5741_elements(138), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2176_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2191_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2206_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2230_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2245_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2271_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2435_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2518_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2543_wire : std_logic_vector(31 downto 0);
    signal LOAD_pad_2114_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2114_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom121_2529_resized : std_logic_vector(13 downto 0);
    signal R_idxprom121_2529_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom126_2554_resized : std_logic_vector(13 downto 0);
    signal R_idxprom126_2554_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2446_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2446_scaled : std_logic_vector(13 downto 0);
    signal add102_2491 : std_logic_vector(31 downto 0);
    signal add112_2506 : std_logic_vector(31 downto 0);
    signal add118_2511 : std_logic_vector(31 downto 0);
    signal add131_2574 : std_logic_vector(31 downto 0);
    signal add139_2594 : std_logic_vector(15 downto 0);
    signal add149_2630 : std_logic_vector(31 downto 0);
    signal add163_2673 : std_logic_vector(31 downto 0);
    signal add64_2386 : std_logic_vector(31 downto 0);
    signal add75_2423 : std_logic_vector(31 downto 0);
    signal add81_2428 : std_logic_vector(31 downto 0);
    signal add93_2486 : std_logic_vector(31 downto 0);
    signal add_2332 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2447_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2447_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2447_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2447_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2447_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2447_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2530_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2530_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2530_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2530_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2530_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2530_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2555_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2555_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2555_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2555_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2555_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2555_root_address : std_logic_vector(13 downto 0);
    signal arrayidx122_2532 : std_logic_vector(31 downto 0);
    signal arrayidx127_2557 : std_logic_vector(31 downto 0);
    signal arrayidx_2449 : std_logic_vector(31 downto 0);
    signal call_2089 : std_logic_vector(15 downto 0);
    signal cmp134_2581 : std_logic_vector(0 downto 0);
    signal cmp150_2635 : std_logic_vector(0 downto 0);
    signal cmp164_2678 : std_logic_vector(0 downto 0);
    signal cmp48_2337 : std_logic_vector(0 downto 0);
    signal cmp55_2356 : std_logic_vector(0 downto 0);
    signal cmp65_2391 : std_logic_vector(0 downto 0);
    signal cmp_2308 : std_logic_vector(0 downto 0);
    signal conv130_2568 : std_logic_vector(31 downto 0);
    signal conv133_2247 : std_logic_vector(31 downto 0);
    signal conv144_2607 : std_logic_vector(31 downto 0);
    signal conv158_2656 : std_logic_vector(31 downto 0);
    signal conv26_2178 : std_logic_vector(31 downto 0);
    signal conv30_2193 : std_logic_vector(31 downto 0);
    signal conv32_2208 : std_logic_vector(31 downto 0);
    signal conv39_2301 : std_logic_vector(31 downto 0);
    signal conv41_2217 : std_logic_vector(31 downto 0);
    signal conv52_2349 : std_logic_vector(31 downto 0);
    signal conv69_2403 : std_logic_vector(31 downto 0);
    signal conv73_2408 : std_logic_vector(31 downto 0);
    signal conv77_2232 : std_logic_vector(31 downto 0);
    signal conv85_2461 : std_logic_vector(31 downto 0);
    signal conv95_2273 : std_logic_vector(31 downto 0);
    signal conv_2112 : std_logic_vector(15 downto 0);
    signal div146_2625 : std_logic_vector(31 downto 0);
    signal div61_2381 : std_logic_vector(31 downto 0);
    signal div_2108 : std_logic_vector(31 downto 0);
    signal iNsTr_11_2323 : std_logic_vector(31 downto 0);
    signal iNsTr_16_2615 : std_logic_vector(31 downto 0);
    signal iNsTr_17_2664 : std_logic_vector(31 downto 0);
    signal iNsTr_19_2371 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2098 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2123 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2135 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2147 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2159 : std_logic_vector(31 downto 0);
    signal idxprom121_2525 : std_logic_vector(63 downto 0);
    signal idxprom126_2550 : std_logic_vector(63 downto 0);
    signal idxprom_2442 : std_logic_vector(63 downto 0);
    signal inc155_2639 : std_logic_vector(15 downto 0);
    signal inc155x_xix_x2_2644 : std_logic_vector(15 downto 0);
    signal inc_2602 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_2686 : std_logic_vector(15 downto 0);
    signal ix_x2_2276 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_2692 : std_logic_vector(15 downto 0);
    signal jx_x1_2282 : std_logic_vector(15 downto 0);
    signal jx_x2_2651 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_2698 : std_logic_vector(15 downto 0);
    signal kx_x1_2289 : std_logic_vector(15 downto 0);
    signal mul101_2481 : std_logic_vector(31 downto 0);
    signal mul111_2496 : std_logic_vector(31 downto 0);
    signal mul117_2501 : std_logic_vector(31 downto 0);
    signal mul33_2213 : std_logic_vector(31 downto 0);
    signal mul74_2413 : std_logic_vector(31 downto 0);
    signal mul80_2418 : std_logic_vector(31 downto 0);
    signal mul92_2471 : std_logic_vector(31 downto 0);
    signal mul_2259 : std_logic_vector(31 downto 0);
    signal ptr_deref_2101_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2101_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2101_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2101_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2101_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2126_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2126_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2126_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2126_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2126_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2138_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2138_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2138_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2138_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2138_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2150_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2150_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2150_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2150_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2150_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2162_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2162_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2162_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2162_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2162_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2326_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2326_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2326_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2326_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2326_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2374_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2374_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2374_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2374_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2374_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2451_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2451_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2451_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2451_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2451_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2451_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2535_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2559_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2559_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2618_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2618_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2618_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2618_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2618_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2667_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2667_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2667_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2667_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2667_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext174_2199 : std_logic_vector(31 downto 0);
    signal sext175_2264 : std_logic_vector(31 downto 0);
    signal sext181_2184 : std_logic_vector(31 downto 0);
    signal sext182_2223 : std_logic_vector(31 downto 0);
    signal sext183_2238 : std_logic_vector(31 downto 0);
    signal sext_2169 : std_logic_vector(31 downto 0);
    signal shl_2253 : std_logic_vector(31 downto 0);
    signal shr120_2520 : std_logic_vector(31 downto 0);
    signal shr125_2545 : std_logic_vector(31 downto 0);
    signal shr_2437 : std_logic_vector(31 downto 0);
    signal sub100_2476 : std_logic_vector(31 downto 0);
    signal sub_2466 : std_logic_vector(31 downto 0);
    signal tmp123_2536 : std_logic_vector(63 downto 0);
    signal tmp145_2619 : std_logic_vector(31 downto 0);
    signal tmp14_2151 : std_logic_vector(31 downto 0);
    signal tmp159_2668 : std_logic_vector(31 downto 0);
    signal tmp17_2163 : std_logic_vector(31 downto 0);
    signal tmp2_2115 : std_logic_vector(7 downto 0);
    signal tmp45_2327 : std_logic_vector(31 downto 0);
    signal tmp5_2127 : std_logic_vector(31 downto 0);
    signal tmp60_2375 : std_logic_vector(31 downto 0);
    signal tmp8_2139 : std_logic_vector(31 downto 0);
    signal tmp_2102 : std_logic_vector(31 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2167_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2172_wire : std_logic_vector(31 downto 0);
    signal type_cast_2175_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2182_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2187_wire : std_logic_vector(31 downto 0);
    signal type_cast_2190_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2202_wire : std_logic_vector(31 downto 0);
    signal type_cast_2205_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2221_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2226_wire : std_logic_vector(31 downto 0);
    signal type_cast_2229_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2236_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2241_wire : std_logic_vector(31 downto 0);
    signal type_cast_2244_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2257_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2267_wire : std_logic_vector(31 downto 0);
    signal type_cast_2270_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2279_wire : std_logic_vector(15 downto 0);
    signal type_cast_2281_wire : std_logic_vector(15 downto 0);
    signal type_cast_2286_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2288_wire : std_logic_vector(15 downto 0);
    signal type_cast_2293_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2295_wire : std_logic_vector(15 downto 0);
    signal type_cast_2299_wire : std_logic_vector(31 downto 0);
    signal type_cast_2304_wire : std_logic_vector(31 downto 0);
    signal type_cast_2306_wire : std_logic_vector(31 downto 0);
    signal type_cast_2347_wire : std_logic_vector(31 downto 0);
    signal type_cast_2352_wire : std_logic_vector(31 downto 0);
    signal type_cast_2354_wire : std_logic_vector(31 downto 0);
    signal type_cast_2379_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2401_wire : std_logic_vector(31 downto 0);
    signal type_cast_2406_wire : std_logic_vector(31 downto 0);
    signal type_cast_2431_wire : std_logic_vector(31 downto 0);
    signal type_cast_2434_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2440_wire : std_logic_vector(63 downto 0);
    signal type_cast_2453_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2459_wire : std_logic_vector(31 downto 0);
    signal type_cast_2514_wire : std_logic_vector(31 downto 0);
    signal type_cast_2517_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2523_wire : std_logic_vector(63 downto 0);
    signal type_cast_2539_wire : std_logic_vector(31 downto 0);
    signal type_cast_2542_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2548_wire : std_logic_vector(63 downto 0);
    signal type_cast_2566_wire : std_logic_vector(31 downto 0);
    signal type_cast_2572_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2577_wire : std_logic_vector(31 downto 0);
    signal type_cast_2579_wire : std_logic_vector(31 downto 0);
    signal type_cast_2592_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2600_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2605_wire : std_logic_vector(31 downto 0);
    signal type_cast_2623_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2648_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2654_wire : std_logic_vector(31 downto 0);
    signal type_cast_2689_wire : std_logic_vector(15 downto 0);
    signal type_cast_2691_wire : std_logic_vector(15 downto 0);
    signal type_cast_2695_wire : std_logic_vector(15 downto 0);
    signal type_cast_2697_wire : std_logic_vector(15 downto 0);
    signal type_cast_2701_wire : std_logic_vector(15 downto 0);
    signal type_cast_2704_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_pad_2114_word_address_0 <= "0";
    array_obj_ref_2447_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2447_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2447_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2447_resized_base_address <= "00000000000000";
    array_obj_ref_2530_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2530_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2530_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2530_resized_base_address <= "00000000000000";
    array_obj_ref_2555_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2555_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2555_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2555_resized_base_address <= "00000000000000";
    iNsTr_11_2323 <= "00000000000000000000000000000011";
    iNsTr_16_2615 <= "00000000000000000000000000000100";
    iNsTr_17_2664 <= "00000000000000000000000000000011";
    iNsTr_19_2371 <= "00000000000000000000000000000100";
    iNsTr_2_2098 <= "00000000000000000000000000000011";
    iNsTr_3_2123 <= "00000000000000000000000000000101";
    iNsTr_4_2135 <= "00000000000000000000000000000100";
    iNsTr_5_2147 <= "00000000000000000000000000000101";
    iNsTr_6_2159 <= "00000000000000000000000000000100";
    ptr_deref_2101_word_offset_0 <= "0000000";
    ptr_deref_2126_word_offset_0 <= "0000000";
    ptr_deref_2138_word_offset_0 <= "0000000";
    ptr_deref_2150_word_offset_0 <= "0000000";
    ptr_deref_2162_word_offset_0 <= "0000000";
    ptr_deref_2326_word_offset_0 <= "0000000";
    ptr_deref_2374_word_offset_0 <= "0000000";
    ptr_deref_2451_word_offset_0 <= "00000000000000";
    ptr_deref_2535_word_offset_0 <= "00000000000000";
    ptr_deref_2559_word_offset_0 <= "00000000000000";
    ptr_deref_2618_word_offset_0 <= "0000000";
    ptr_deref_2667_word_offset_0 <= "0000000";
    type_cast_2106_wire_constant <= "00000000000000000000000000000001";
    type_cast_2167_wire_constant <= "00000000000000000000000000010000";
    type_cast_2175_wire_constant <= "00000000000000000000000000010000";
    type_cast_2182_wire_constant <= "00000000000000000000000000010000";
    type_cast_2190_wire_constant <= "00000000000000000000000000010000";
    type_cast_2197_wire_constant <= "00000000000000000000000000010000";
    type_cast_2205_wire_constant <= "00000000000000000000000000010000";
    type_cast_2221_wire_constant <= "00000000000000000000000000010000";
    type_cast_2229_wire_constant <= "00000000000000000000000000010000";
    type_cast_2236_wire_constant <= "00000000000000000000000000010000";
    type_cast_2244_wire_constant <= "00000000000000000000000000010000";
    type_cast_2251_wire_constant <= "00000000000000000000000000000001";
    type_cast_2257_wire_constant <= "00000000000000000000000000010000";
    type_cast_2270_wire_constant <= "00000000000000000000000000010000";
    type_cast_2286_wire_constant <= "0000000000000000";
    type_cast_2293_wire_constant <= "0000000000000000";
    type_cast_2379_wire_constant <= "00000000000000000000000000000001";
    type_cast_2434_wire_constant <= "00000000000000000000000000000010";
    type_cast_2453_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2517_wire_constant <= "00000000000000000000000000000010";
    type_cast_2542_wire_constant <= "00000000000000000000000000000010";
    type_cast_2572_wire_constant <= "00000000000000000000000000000100";
    type_cast_2592_wire_constant <= "0000000000000100";
    type_cast_2600_wire_constant <= "0000000000000001";
    type_cast_2623_wire_constant <= "00000000000000000000000000000001";
    type_cast_2648_wire_constant <= "0000000000000000";
    type_cast_2704_wire_constant <= "0000000000000000";
    phi_stmt_2276: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2279_wire & type_cast_2281_wire;
      req <= phi_stmt_2276_req_0 & phi_stmt_2276_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2276",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2276_ack_0,
          idata => idata,
          odata => ix_x2_2276,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2276
    phi_stmt_2282: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2286_wire_constant & type_cast_2288_wire;
      req <= phi_stmt_2282_req_0 & phi_stmt_2282_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2282",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2282_ack_0,
          idata => idata,
          odata => jx_x1_2282,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2282
    phi_stmt_2289: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2293_wire_constant & type_cast_2295_wire;
      req <= phi_stmt_2289_req_0 & phi_stmt_2289_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2289",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2289_ack_0,
          idata => idata,
          odata => kx_x1_2289,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2289
    phi_stmt_2686: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2689_wire & type_cast_2691_wire;
      req <= phi_stmt_2686_req_0 & phi_stmt_2686_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2686",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2686_ack_0,
          idata => idata,
          odata => ix_x1x_xph_2686,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2686
    phi_stmt_2692: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2695_wire & type_cast_2697_wire;
      req <= phi_stmt_2692_req_0 & phi_stmt_2692_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2692",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2692_ack_0,
          idata => idata,
          odata => jx_x0x_xph_2692,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2692
    phi_stmt_2698: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2701_wire & type_cast_2704_wire_constant;
      req <= phi_stmt_2698_req_0 & phi_stmt_2698_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2698",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2698_ack_0,
          idata => idata,
          odata => kx_x0x_xph_2698,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2698
    -- flow-through select operator MUX_2650_inst
    jx_x2_2651 <= type_cast_2648_wire_constant when (cmp150_2635(0) /=  '0') else inc_2602;
    addr_of_2448_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2448_final_reg_req_0;
      addr_of_2448_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2448_final_reg_req_1;
      addr_of_2448_final_reg_ack_1<= rack(0);
      addr_of_2448_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2448_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2447_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2531_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2531_final_reg_req_0;
      addr_of_2531_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2531_final_reg_req_1;
      addr_of_2531_final_reg_ack_1<= rack(0);
      addr_of_2531_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2531_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2530_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx122_2532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2556_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2556_final_reg_req_0;
      addr_of_2556_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2556_final_reg_req_1;
      addr_of_2556_final_reg_ack_1<= rack(0);
      addr_of_2556_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2556_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2555_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx127_2557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2111_inst_req_0;
      type_cast_2111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2111_inst_req_1;
      type_cast_2111_inst_ack_1<= rack(0);
      type_cast_2111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2172_inst
    process(sext_2169) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2169(31 downto 0);
      type_cast_2172_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2177_inst
    process(ASHR_i32_i32_2176_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2176_wire(31 downto 0);
      conv26_2178 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2187_inst
    process(sext181_2184) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext181_2184(31 downto 0);
      type_cast_2187_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2192_inst
    process(ASHR_i32_i32_2191_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2191_wire(31 downto 0);
      conv30_2193 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2202_inst
    process(sext174_2199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext174_2199(31 downto 0);
      type_cast_2202_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2207_inst
    process(ASHR_i32_i32_2206_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2206_wire(31 downto 0);
      conv32_2208 <= tmp_var; -- 
    end process;
    type_cast_2216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2216_inst_req_0;
      type_cast_2216_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2216_inst_req_1;
      type_cast_2216_inst_ack_1<= rack(0);
      type_cast_2216_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2216_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp2_2115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_2217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2226_inst
    process(sext182_2223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext182_2223(31 downto 0);
      type_cast_2226_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2231_inst
    process(ASHR_i32_i32_2230_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2230_wire(31 downto 0);
      conv77_2232 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2241_inst
    process(sext183_2238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext183_2238(31 downto 0);
      type_cast_2241_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2246_inst
    process(ASHR_i32_i32_2245_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2245_wire(31 downto 0);
      conv133_2247 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2267_inst
    process(sext175_2264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext175_2264(31 downto 0);
      type_cast_2267_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2272_inst
    process(ASHR_i32_i32_2271_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2271_wire(31 downto 0);
      conv95_2273 <= tmp_var; -- 
    end process;
    type_cast_2279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2279_inst_req_0;
      type_cast_2279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2279_inst_req_1;
      type_cast_2279_inst_ack_1<= rack(0);
      type_cast_2279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2279_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2281_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2281_inst_req_0;
      type_cast_2281_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2281_inst_req_1;
      type_cast_2281_inst_ack_1<= rack(0);
      type_cast_2281_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2281_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_2686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2281_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2288_inst_req_0;
      type_cast_2288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2288_inst_req_1;
      type_cast_2288_inst_ack_1<= rack(0);
      type_cast_2288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_2692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2288_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2295_inst_req_0;
      type_cast_2295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2295_inst_req_1;
      type_cast_2295_inst_ack_1<= rack(0);
      type_cast_2295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_2698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2295_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2300_inst_req_0;
      type_cast_2300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2300_inst_req_1;
      type_cast_2300_inst_ack_1<= rack(0);
      type_cast_2300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2299_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_2301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2304_inst
    process(conv39_2301) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv39_2301(31 downto 0);
      type_cast_2304_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2306_inst
    process(conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv41_2217(31 downto 0);
      type_cast_2306_wire <= tmp_var; -- 
    end process;
    type_cast_2348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2348_inst_req_0;
      type_cast_2348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2348_inst_req_1;
      type_cast_2348_inst_ack_1<= rack(0);
      type_cast_2348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2347_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_2349,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2352_inst
    process(conv52_2349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv52_2349(31 downto 0);
      type_cast_2352_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2354_inst
    process(conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv41_2217(31 downto 0);
      type_cast_2354_wire <= tmp_var; -- 
    end process;
    type_cast_2402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2402_inst_req_0;
      type_cast_2402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2402_inst_req_1;
      type_cast_2402_inst_ack_1<= rack(0);
      type_cast_2402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2401_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_2403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2407_inst_req_0;
      type_cast_2407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2407_inst_req_1;
      type_cast_2407_inst_ack_1<= rack(0);
      type_cast_2407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2406_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2408,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2431_inst
    process(add81_2428) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add81_2428(31 downto 0);
      type_cast_2431_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2436_inst
    process(ASHR_i32_i32_2435_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2435_wire(31 downto 0);
      shr_2437 <= tmp_var; -- 
    end process;
    type_cast_2441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2441_inst_req_0;
      type_cast_2441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2441_inst_req_1;
      type_cast_2441_inst_ack_1<= rack(0);
      type_cast_2441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2440_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2460_inst_req_0;
      type_cast_2460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2460_inst_req_1;
      type_cast_2460_inst_ack_1<= rack(0);
      type_cast_2460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2459_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2461,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2514_inst
    process(add102_2491) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add102_2491(31 downto 0);
      type_cast_2514_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2519_inst
    process(ASHR_i32_i32_2518_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2518_wire(31 downto 0);
      shr120_2520 <= tmp_var; -- 
    end process;
    type_cast_2524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2524_inst_req_0;
      type_cast_2524_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2524_inst_req_1;
      type_cast_2524_inst_ack_1<= rack(0);
      type_cast_2524_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2524_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2523_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom121_2525,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2539_inst
    process(add118_2511) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add118_2511(31 downto 0);
      type_cast_2539_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2544_inst
    process(ASHR_i32_i32_2543_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2543_wire(31 downto 0);
      shr125_2545 <= tmp_var; -- 
    end process;
    type_cast_2549_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2549_inst_req_0;
      type_cast_2549_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2549_inst_req_1;
      type_cast_2549_inst_ack_1<= rack(0);
      type_cast_2549_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2549_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2548_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom126_2550,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2567_inst_req_0;
      type_cast_2567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2567_inst_req_1;
      type_cast_2567_inst_ack_1<= rack(0);
      type_cast_2567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2566_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_2568,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2577_inst
    process(add131_2574) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add131_2574(31 downto 0);
      type_cast_2577_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2579_inst
    process(conv133_2247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv133_2247(31 downto 0);
      type_cast_2579_wire <= tmp_var; -- 
    end process;
    type_cast_2606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2606_inst_req_0;
      type_cast_2606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2606_inst_req_1;
      type_cast_2606_inst_ack_1<= rack(0);
      type_cast_2606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2605_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_2607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2638_inst_req_0;
      type_cast_2638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2638_inst_req_1;
      type_cast_2638_inst_ack_1<= rack(0);
      type_cast_2638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp150_2635,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc155_2639,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2655_inst_req_0;
      type_cast_2655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2655_inst_req_1;
      type_cast_2655_inst_ack_1<= rack(0);
      type_cast_2655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2654_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_2656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2689_inst_req_0;
      type_cast_2689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2689_inst_req_1;
      type_cast_2689_inst_ack_1<= rack(0);
      type_cast_2689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_2276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2689_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2691_inst_req_0;
      type_cast_2691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2691_inst_req_1;
      type_cast_2691_inst_ack_1<= rack(0);
      type_cast_2691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc155x_xix_x2_2644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2691_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2695_inst_req_0;
      type_cast_2695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2695_inst_req_1;
      type_cast_2695_inst_ack_1<= rack(0);
      type_cast_2695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_2282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2695_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2697_inst_req_0;
      type_cast_2697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2697_inst_req_1;
      type_cast_2697_inst_ack_1<= rack(0);
      type_cast_2697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_2651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2697_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2701_inst_req_0;
      type_cast_2701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2701_inst_req_1;
      type_cast_2701_inst_ack_1<= rack(0);
      type_cast_2701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add139_2594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2701_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_pad_2114_gather_scatter
    process(LOAD_pad_2114_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2114_data_0;
      ov(7 downto 0) := iv;
      tmp2_2115 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2447_index_1_rename
    process(R_idxprom_2446_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2446_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2446_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2447_index_1_resize
    process(idxprom_2442) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2442;
      ov := iv(13 downto 0);
      R_idxprom_2446_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2447_root_address_inst
    process(array_obj_ref_2447_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2447_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2447_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2530_index_1_rename
    process(R_idxprom121_2529_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom121_2529_resized;
      ov(13 downto 0) := iv;
      R_idxprom121_2529_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2530_index_1_resize
    process(idxprom121_2525) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom121_2525;
      ov := iv(13 downto 0);
      R_idxprom121_2529_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2530_root_address_inst
    process(array_obj_ref_2530_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2530_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2530_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2555_index_1_rename
    process(R_idxprom126_2554_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom126_2554_resized;
      ov(13 downto 0) := iv;
      R_idxprom126_2554_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2555_index_1_resize
    process(idxprom126_2550) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom126_2550;
      ov := iv(13 downto 0);
      R_idxprom126_2554_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2555_root_address_inst
    process(array_obj_ref_2555_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2555_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2555_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_addr_0
    process(ptr_deref_2101_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2101_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_base_resize
    process(iNsTr_2_2098) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2098;
      ov := iv(6 downto 0);
      ptr_deref_2101_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_gather_scatter
    process(ptr_deref_2101_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_data_0;
      ov(31 downto 0) := iv;
      tmp_2102 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_root_address_inst
    process(ptr_deref_2101_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2101_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2126_addr_0
    process(ptr_deref_2126_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2126_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2126_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2126_base_resize
    process(iNsTr_3_2123) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2123;
      ov := iv(6 downto 0);
      ptr_deref_2126_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2126_gather_scatter
    process(ptr_deref_2126_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2126_data_0;
      ov(31 downto 0) := iv;
      tmp5_2127 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2126_root_address_inst
    process(ptr_deref_2126_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2126_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2126_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2138_addr_0
    process(ptr_deref_2138_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2138_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2138_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2138_base_resize
    process(iNsTr_4_2135) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2135;
      ov := iv(6 downto 0);
      ptr_deref_2138_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2138_gather_scatter
    process(ptr_deref_2138_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2138_data_0;
      ov(31 downto 0) := iv;
      tmp8_2139 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2138_root_address_inst
    process(ptr_deref_2138_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2138_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2138_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_addr_0
    process(ptr_deref_2150_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2150_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2150_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_base_resize
    process(iNsTr_5_2147) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2147;
      ov := iv(6 downto 0);
      ptr_deref_2150_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_gather_scatter
    process(ptr_deref_2150_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2150_data_0;
      ov(31 downto 0) := iv;
      tmp14_2151 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_root_address_inst
    process(ptr_deref_2150_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2150_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2150_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2162_addr_0
    process(ptr_deref_2162_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2162_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2162_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2162_base_resize
    process(iNsTr_6_2159) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2159;
      ov := iv(6 downto 0);
      ptr_deref_2162_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2162_gather_scatter
    process(ptr_deref_2162_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2162_data_0;
      ov(31 downto 0) := iv;
      tmp17_2163 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2162_root_address_inst
    process(ptr_deref_2162_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2162_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2162_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2326_addr_0
    process(ptr_deref_2326_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2326_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2326_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2326_base_resize
    process(iNsTr_11_2323) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_11_2323;
      ov := iv(6 downto 0);
      ptr_deref_2326_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2326_gather_scatter
    process(ptr_deref_2326_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2326_data_0;
      ov(31 downto 0) := iv;
      tmp45_2327 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2326_root_address_inst
    process(ptr_deref_2326_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2326_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2326_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2374_addr_0
    process(ptr_deref_2374_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2374_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2374_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2374_base_resize
    process(iNsTr_19_2371) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_19_2371;
      ov := iv(6 downto 0);
      ptr_deref_2374_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2374_gather_scatter
    process(ptr_deref_2374_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2374_data_0;
      ov(31 downto 0) := iv;
      tmp60_2375 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2374_root_address_inst
    process(ptr_deref_2374_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2374_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2374_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_addr_0
    process(ptr_deref_2451_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2451_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2451_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_base_resize
    process(arrayidx_2449) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2449;
      ov := iv(13 downto 0);
      ptr_deref_2451_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_gather_scatter
    process(type_cast_2453_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2453_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2451_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_root_address_inst
    process(ptr_deref_2451_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2451_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2451_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_addr_0
    process(ptr_deref_2535_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2535_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2535_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_base_resize
    process(arrayidx122_2532) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx122_2532;
      ov := iv(13 downto 0);
      ptr_deref_2535_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_gather_scatter
    process(ptr_deref_2535_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2535_data_0;
      ov(63 downto 0) := iv;
      tmp123_2536 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_root_address_inst
    process(ptr_deref_2535_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2535_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2535_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_addr_0
    process(ptr_deref_2559_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2559_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2559_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_base_resize
    process(arrayidx127_2557) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx127_2557;
      ov := iv(13 downto 0);
      ptr_deref_2559_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_gather_scatter
    process(tmp123_2536) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp123_2536;
      ov(63 downto 0) := iv;
      ptr_deref_2559_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_root_address_inst
    process(ptr_deref_2559_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2559_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2559_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2618_addr_0
    process(ptr_deref_2618_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2618_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2618_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2618_base_resize
    process(iNsTr_16_2615) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_16_2615;
      ov := iv(6 downto 0);
      ptr_deref_2618_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2618_gather_scatter
    process(ptr_deref_2618_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2618_data_0;
      ov(31 downto 0) := iv;
      tmp145_2619 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2618_root_address_inst
    process(ptr_deref_2618_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2618_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2618_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2667_addr_0
    process(ptr_deref_2667_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2667_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2667_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2667_base_resize
    process(iNsTr_17_2664) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_2664;
      ov := iv(6 downto 0);
      ptr_deref_2667_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2667_gather_scatter
    process(ptr_deref_2667_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2667_data_0;
      ov(31 downto 0) := iv;
      tmp159_2668 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2667_root_address_inst
    process(ptr_deref_2667_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2667_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2667_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_2309_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2308;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2309_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2309_branch_req_0,
          ack0 => if_stmt_2309_branch_ack_0,
          ack1 => if_stmt_2309_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2338_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp48_2337;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2338_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2338_branch_req_0,
          ack0 => if_stmt_2338_branch_ack_0,
          ack1 => if_stmt_2338_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2357_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp55_2356;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2357_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2357_branch_req_0,
          ack0 => if_stmt_2357_branch_ack_0,
          ack1 => if_stmt_2357_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2392_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp65_2391;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2392_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2392_branch_req_0,
          ack0 => if_stmt_2392_branch_ack_0,
          ack1 => if_stmt_2392_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2582_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp134_2581;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2582_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2582_branch_req_0,
          ack0 => if_stmt_2582_branch_ack_0,
          ack1 => if_stmt_2582_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2679_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp164_2678;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2679_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2679_branch_req_0,
          ack0 => if_stmt_2679_branch_ack_0,
          ack1 => if_stmt_2679_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2593_inst
    process(kx_x1_2289) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_2289, type_cast_2592_wire_constant, tmp_var);
      add139_2594 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2601_inst
    process(jx_x1_2282) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_2282, type_cast_2600_wire_constant, tmp_var);
      inc_2602 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2643_inst
    process(inc155_2639, ix_x2_2276) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc155_2639, ix_x2_2276, tmp_var);
      inc155x_xix_x2_2644 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2331_inst
    process(tmp45_2327, conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp45_2327, conv41_2217, tmp_var);
      add_2332 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2385_inst
    process(div61_2381, conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div61_2381, conv41_2217, tmp_var);
      add64_2386 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2422_inst
    process(mul74_2413, mul80_2418) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_2413, mul80_2418, tmp_var);
      add75_2423 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2427_inst
    process(add75_2423, conv69_2403) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add75_2423, conv69_2403, tmp_var);
      add81_2428 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2485_inst
    process(conv85_2461, mul101_2481) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_2461, mul101_2481, tmp_var);
      add93_2486 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2490_inst
    process(add93_2486, mul92_2471) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add93_2486, mul92_2471, tmp_var);
      add102_2491 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2505_inst
    process(mul111_2496, mul117_2501) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul111_2496, mul117_2501, tmp_var);
      add112_2506 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2510_inst
    process(add112_2506, conv85_2461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add112_2506, conv85_2461, tmp_var);
      add118_2511 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2573_inst
    process(conv130_2568) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv130_2568, type_cast_2572_wire_constant, tmp_var);
      add131_2574 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2629_inst
    process(div146_2625, shl_2253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div146_2625, shl_2253, tmp_var);
      add149_2630 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2672_inst
    process(tmp159_2668, shl_2253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp159_2668, shl_2253, tmp_var);
      add163_2673 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2176_inst
    process(type_cast_2172_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2172_wire, type_cast_2175_wire_constant, tmp_var);
      ASHR_i32_i32_2176_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2191_inst
    process(type_cast_2187_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2187_wire, type_cast_2190_wire_constant, tmp_var);
      ASHR_i32_i32_2191_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2206_inst
    process(type_cast_2202_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2202_wire, type_cast_2205_wire_constant, tmp_var);
      ASHR_i32_i32_2206_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2230_inst
    process(type_cast_2226_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2226_wire, type_cast_2229_wire_constant, tmp_var);
      ASHR_i32_i32_2230_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2245_inst
    process(type_cast_2241_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2241_wire, type_cast_2244_wire_constant, tmp_var);
      ASHR_i32_i32_2245_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2271_inst
    process(type_cast_2267_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2267_wire, type_cast_2270_wire_constant, tmp_var);
      ASHR_i32_i32_2271_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2435_inst
    process(type_cast_2431_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2431_wire, type_cast_2434_wire_constant, tmp_var);
      ASHR_i32_i32_2435_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2518_inst
    process(type_cast_2514_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2514_wire, type_cast_2517_wire_constant, tmp_var);
      ASHR_i32_i32_2518_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2543_inst
    process(type_cast_2539_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2539_wire, type_cast_2542_wire_constant, tmp_var);
      ASHR_i32_i32_2543_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2634_inst
    process(conv144_2607, add149_2630) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv144_2607, add149_2630, tmp_var);
      cmp150_2635 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2677_inst
    process(conv158_2656, add163_2673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv158_2656, add163_2673, tmp_var);
      cmp164_2678 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2107_inst
    process(tmp_2102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2102, type_cast_2106_wire_constant, tmp_var);
      div_2108 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2380_inst
    process(tmp60_2375) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp60_2375, type_cast_2379_wire_constant, tmp_var);
      div61_2381 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2624_inst
    process(tmp145_2619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp145_2619, type_cast_2623_wire_constant, tmp_var);
      div146_2625 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2212_inst
    process(conv32_2208, conv30_2193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv32_2208, conv30_2193, tmp_var);
      mul33_2213 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2263_inst
    process(mul_2259, conv26_2178) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_2259, conv26_2178, tmp_var);
      sext175_2264 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2412_inst
    process(conv73_2408, conv30_2193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv73_2408, conv30_2193, tmp_var);
      mul74_2413 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2417_inst
    process(conv39_2301, conv77_2232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv39_2301, conv77_2232, tmp_var);
      mul80_2418 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2470_inst
    process(sub_2466, conv133_2247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_2466, conv133_2247, tmp_var);
      mul92_2471 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2480_inst
    process(sub100_2476, conv95_2273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub100_2476, conv95_2273, tmp_var);
      mul101_2481 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2495_inst
    process(conv52_2349, conv30_2193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv52_2349, conv30_2193, tmp_var);
      mul111_2496 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2500_inst
    process(conv39_2301, conv77_2232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv39_2301, conv77_2232, tmp_var);
      mul117_2501 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2168_inst
    process(tmp8_2139) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp8_2139, type_cast_2167_wire_constant, tmp_var);
      sext_2169 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2183_inst
    process(tmp14_2151) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp14_2151, type_cast_2182_wire_constant, tmp_var);
      sext181_2184 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2198_inst
    process(tmp17_2163) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp17_2163, type_cast_2197_wire_constant, tmp_var);
      sext174_2199 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2222_inst
    process(mul33_2213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul33_2213, type_cast_2221_wire_constant, tmp_var);
      sext182_2223 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2237_inst
    process(tmp5_2127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp5_2127, type_cast_2236_wire_constant, tmp_var);
      sext183_2238 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2252_inst
    process(conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv41_2217, type_cast_2251_wire_constant, tmp_var);
      shl_2253 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2258_inst
    process(tmp5_2127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp5_2127, type_cast_2257_wire_constant, tmp_var);
      mul_2259 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2307_inst
    process(type_cast_2304_wire, type_cast_2306_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2304_wire, type_cast_2306_wire, tmp_var);
      cmp_2308 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2355_inst
    process(type_cast_2352_wire, type_cast_2354_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2352_wire, type_cast_2354_wire, tmp_var);
      cmp55_2356 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2580_inst
    process(type_cast_2577_wire, type_cast_2579_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2577_wire, type_cast_2579_wire, tmp_var);
      cmp134_2581 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2465_inst
    process(conv52_2349, conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv52_2349, conv41_2217, tmp_var);
      sub_2466 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2475_inst
    process(conv39_2301, conv41_2217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv39_2301, conv41_2217, tmp_var);
      sub100_2476 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2336_inst
    process(conv39_2301, add_2332) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv39_2301, add_2332, tmp_var);
      cmp48_2337 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2390_inst
    process(conv52_2349, add64_2386) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv52_2349, add64_2386, tmp_var);
      cmp65_2391 <= tmp_var; --
    end process;
    -- shared split operator group (50) : array_obj_ref_2447_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2446_scaled;
      array_obj_ref_2447_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2447_index_offset_req_0;
      array_obj_ref_2447_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2447_index_offset_req_1;
      array_obj_ref_2447_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : array_obj_ref_2530_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom121_2529_scaled;
      array_obj_ref_2530_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2530_index_offset_req_0;
      array_obj_ref_2530_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2530_index_offset_req_1;
      array_obj_ref_2530_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : array_obj_ref_2555_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom126_2554_scaled;
      array_obj_ref_2555_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2555_index_offset_req_0;
      array_obj_ref_2555_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2555_index_offset_req_1;
      array_obj_ref_2555_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- unary operator type_cast_2299_inst
    process(ix_x2_2276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_2276, tmp_var);
      type_cast_2299_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2347_inst
    process(jx_x1_2282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2282, tmp_var);
      type_cast_2347_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2401_inst
    process(kx_x1_2289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2289, tmp_var);
      type_cast_2401_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2406_inst
    process(jx_x1_2282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2282, tmp_var);
      type_cast_2406_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2440_inst
    process(shr_2437) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2437, tmp_var);
      type_cast_2440_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2459_inst
    process(kx_x1_2289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2289, tmp_var);
      type_cast_2459_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2523_inst
    process(shr120_2520) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr120_2520, tmp_var);
      type_cast_2523_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2548_inst
    process(shr125_2545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr125_2545, tmp_var);
      type_cast_2548_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2566_inst
    process(kx_x1_2289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2289, tmp_var);
      type_cast_2566_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2605_inst
    process(inc_2602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2602, tmp_var);
      type_cast_2605_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2654_inst
    process(inc155x_xix_x2_2644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc155x_xix_x2_2644, tmp_var);
      type_cast_2654_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_pad_2114_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_pad_2114_load_0_req_0;
      LOAD_pad_2114_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_pad_2114_load_0_req_1;
      LOAD_pad_2114_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_2114_word_address_0;
      LOAD_pad_2114_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(0 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2374_load_0 ptr_deref_2326_load_0 ptr_deref_2667_load_0 ptr_deref_2618_load_0 ptr_deref_2101_load_0 ptr_deref_2126_load_0 ptr_deref_2138_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(48 downto 0);
      signal data_out: std_logic_vector(223 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= ptr_deref_2374_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_2326_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_2667_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2618_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_2101_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2126_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2138_load_0_req_0;
      ptr_deref_2374_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_2326_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_2667_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2618_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_2101_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2126_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2138_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= ptr_deref_2374_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_2326_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_2667_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2618_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_2101_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2126_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2138_load_0_req_1;
      ptr_deref_2374_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_2326_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_2667_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2618_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_2101_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2126_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2138_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2374_word_address_0 & ptr_deref_2326_word_address_0 & ptr_deref_2667_word_address_0 & ptr_deref_2618_word_address_0 & ptr_deref_2101_word_address_0 & ptr_deref_2126_word_address_0 & ptr_deref_2138_word_address_0;
      ptr_deref_2374_data_0 <= data_out(223 downto 192);
      ptr_deref_2326_data_0 <= data_out(191 downto 160);
      ptr_deref_2667_data_0 <= data_out(159 downto 128);
      ptr_deref_2618_data_0 <= data_out(127 downto 96);
      ptr_deref_2101_data_0 <= data_out(95 downto 64);
      ptr_deref_2126_data_0 <= data_out(63 downto 32);
      ptr_deref_2138_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 7,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 7,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2162_load_0 ptr_deref_2150_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2162_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2150_load_0_req_0;
      ptr_deref_2162_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2150_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2162_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2150_load_0_req_1;
      ptr_deref_2162_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2150_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2162_word_address_0 & ptr_deref_2150_word_address_0;
      ptr_deref_2162_data_0 <= data_out(63 downto 32);
      ptr_deref_2150_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(6 downto 0),
          mtag => memory_space_4_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2535_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2535_load_0_req_0;
      ptr_deref_2535_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2535_load_0_req_1;
      ptr_deref_2535_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2535_word_address_0;
      ptr_deref_2535_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_2451_store_0 ptr_deref_2559_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2451_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2559_store_0_req_0;
      ptr_deref_2451_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2559_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2451_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2559_store_0_req_1;
      ptr_deref_2451_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2559_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2451_word_address_0 & ptr_deref_2559_word_address_0;
      data_in <= ptr_deref_2451_data_0 & ptr_deref_2559_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_starting_2088_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_starting_2088_inst_req_0;
      RPIPE_Block2_starting_2088_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_starting_2088_inst_req_1;
      RPIPE_Block2_starting_2088_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2089 <= data_out(15 downto 0);
      Block2_starting_read_0_gI: SplitGuardInterface generic map(name => "Block2_starting_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block2_starting_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_starting_pipe_read_req(0),
          oack => Block2_starting_pipe_read_ack(0),
          odata => Block2_starting_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_complete_2709_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_complete_2709_inst_req_0;
      WPIPE_Block2_complete_2709_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_complete_2709_inst_req_1;
      WPIPE_Block2_complete_2709_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2089;
      Block2_complete_write_0_gI: SplitGuardInterface generic map(name => "Block2_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_complete", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_complete_pipe_write_req(0),
          oack => Block2_complete_pipe_write_ack(0),
          odata => Block2_complete_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_C_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block3_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_D;
architecture zeropad3D_D_arch of zeropad3D_D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_D_CP_7327_start: Boolean;
  signal zeropad3D_D_CP_7327_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2764_inst_req_0 : boolean;
  signal type_cast_2764_inst_ack_0 : boolean;
  signal LOAD_pad_2767_load_0_ack_1 : boolean;
  signal type_cast_2764_inst_req_1 : boolean;
  signal type_cast_2764_inst_ack_1 : boolean;
  signal ptr_deref_2754_load_0_req_1 : boolean;
  signal ptr_deref_2754_load_0_ack_1 : boolean;
  signal ptr_deref_2754_load_0_req_0 : boolean;
  signal ptr_deref_2732_load_0_req_1 : boolean;
  signal ptr_deref_2732_load_0_ack_1 : boolean;
  signal ptr_deref_2732_load_0_ack_0 : boolean;
  signal LOAD_pad_2767_load_0_req_0 : boolean;
  signal LOAD_pad_2767_load_0_ack_0 : boolean;
  signal LOAD_pad_2767_load_0_req_1 : boolean;
  signal type_cast_2742_inst_ack_1 : boolean;
  signal type_cast_2742_inst_req_0 : boolean;
  signal type_cast_2742_inst_req_1 : boolean;
  signal type_cast_2742_inst_ack_0 : boolean;
  signal ptr_deref_2779_load_0_req_0 : boolean;
  signal ptr_deref_2732_load_0_req_0 : boolean;
  signal ptr_deref_2754_load_0_ack_0 : boolean;
  signal phi_stmt_2923_req_0 : boolean;
  signal ptr_deref_3294_load_0_req_1 : boolean;
  signal phi_stmt_2929_req_0 : boolean;
  signal type_cast_2922_inst_ack_0 : boolean;
  signal type_cast_3266_inst_req_0 : boolean;
  signal type_cast_2926_inst_req_1 : boolean;
  signal ptr_deref_3193_store_0_req_1 : boolean;
  signal type_cast_2928_inst_req_0 : boolean;
  signal ptr_deref_3193_store_0_req_0 : boolean;
  signal type_cast_2922_inst_req_0 : boolean;
  signal type_cast_2926_inst_ack_1 : boolean;
  signal type_cast_3266_inst_ack_0 : boolean;
  signal ptr_deref_3193_store_0_ack_1 : boolean;
  signal ptr_deref_3294_load_0_req_0 : boolean;
  signal type_cast_2928_inst_req_1 : boolean;
  signal type_cast_2928_inst_ack_1 : boolean;
  signal ptr_deref_3294_load_0_ack_1 : boolean;
  signal type_cast_2935_inst_req_1 : boolean;
  signal type_cast_2935_inst_ack_1 : boolean;
  signal phi_stmt_2929_req_1 : boolean;
  signal phi_stmt_2917_ack_0 : boolean;
  signal phi_stmt_2923_ack_0 : boolean;
  signal phi_stmt_2929_ack_0 : boolean;
  signal type_cast_2926_inst_ack_0 : boolean;
  signal type_cast_3266_inst_req_1 : boolean;
  signal type_cast_3266_inst_ack_1 : boolean;
  signal ptr_deref_3294_load_0_ack_0 : boolean;
  signal type_cast_2920_inst_req_0 : boolean;
  signal ptr_deref_3193_store_0_ack_0 : boolean;
  signal type_cast_2926_inst_req_0 : boolean;
  signal phi_stmt_2923_req_1 : boolean;
  signal type_cast_2928_inst_ack_0 : boolean;
  signal type_cast_3240_inst_req_0 : boolean;
  signal type_cast_2920_inst_ack_0 : boolean;
  signal type_cast_2935_inst_req_0 : boolean;
  signal type_cast_2935_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2719_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2719_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2719_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2719_inst_ack_1 : boolean;
  signal ptr_deref_2779_load_0_ack_0 : boolean;
  signal ptr_deref_2779_load_0_req_1 : boolean;
  signal ptr_deref_2779_load_0_ack_1 : boolean;
  signal ptr_deref_2791_load_0_req_0 : boolean;
  signal ptr_deref_2791_load_0_ack_0 : boolean;
  signal ptr_deref_2791_load_0_req_1 : boolean;
  signal ptr_deref_2791_load_0_ack_1 : boolean;
  signal ptr_deref_2803_load_0_req_0 : boolean;
  signal ptr_deref_2803_load_0_ack_0 : boolean;
  signal ptr_deref_2803_load_0_req_1 : boolean;
  signal ptr_deref_2803_load_0_ack_1 : boolean;
  signal type_cast_2857_inst_req_0 : boolean;
  signal type_cast_2857_inst_ack_0 : boolean;
  signal type_cast_2857_inst_req_1 : boolean;
  signal type_cast_2857_inst_ack_1 : boolean;
  signal type_cast_2940_inst_req_0 : boolean;
  signal type_cast_2940_inst_ack_0 : boolean;
  signal type_cast_2940_inst_req_1 : boolean;
  signal type_cast_2940_inst_ack_1 : boolean;
  signal if_stmt_2949_branch_req_0 : boolean;
  signal if_stmt_2949_branch_ack_1 : boolean;
  signal if_stmt_2949_branch_ack_0 : boolean;
  signal ptr_deref_2966_load_0_req_0 : boolean;
  signal ptr_deref_2966_load_0_ack_0 : boolean;
  signal ptr_deref_2966_load_0_req_1 : boolean;
  signal ptr_deref_2966_load_0_ack_1 : boolean;
  signal if_stmt_2978_branch_req_0 : boolean;
  signal if_stmt_2978_branch_ack_1 : boolean;
  signal if_stmt_2978_branch_ack_0 : boolean;
  signal type_cast_2988_inst_req_0 : boolean;
  signal type_cast_2988_inst_ack_0 : boolean;
  signal type_cast_2988_inst_req_1 : boolean;
  signal type_cast_2988_inst_ack_1 : boolean;
  signal if_stmt_2997_branch_req_0 : boolean;
  signal if_stmt_2997_branch_ack_1 : boolean;
  signal if_stmt_2997_branch_ack_0 : boolean;
  signal ptr_deref_3014_load_0_req_0 : boolean;
  signal ptr_deref_3014_load_0_ack_0 : boolean;
  signal ptr_deref_3014_load_0_req_1 : boolean;
  signal ptr_deref_3014_load_0_ack_1 : boolean;
  signal if_stmt_3026_branch_req_0 : boolean;
  signal if_stmt_3026_branch_ack_1 : boolean;
  signal if_stmt_3026_branch_ack_0 : boolean;
  signal type_cast_3036_inst_req_0 : boolean;
  signal type_cast_3036_inst_ack_0 : boolean;
  signal type_cast_3036_inst_req_1 : boolean;
  signal type_cast_3036_inst_ack_1 : boolean;
  signal type_cast_3041_inst_req_0 : boolean;
  signal type_cast_3041_inst_ack_0 : boolean;
  signal if_stmt_3306_branch_ack_0 : boolean;
  signal type_cast_3041_inst_req_1 : boolean;
  signal type_cast_3041_inst_ack_1 : boolean;
  signal ptr_deref_3252_load_0_ack_1 : boolean;
  signal type_cast_3075_inst_req_0 : boolean;
  signal ptr_deref_3252_load_0_req_1 : boolean;
  signal type_cast_3075_inst_ack_0 : boolean;
  signal if_stmt_3306_branch_ack_1 : boolean;
  signal type_cast_3075_inst_req_1 : boolean;
  signal type_cast_3075_inst_ack_1 : boolean;
  signal phi_stmt_2917_req_1 : boolean;
  signal if_stmt_3216_branch_ack_0 : boolean;
  signal type_cast_3240_inst_ack_1 : boolean;
  signal array_obj_ref_3081_index_offset_req_0 : boolean;
  signal array_obj_ref_3081_index_offset_ack_0 : boolean;
  signal array_obj_ref_3081_index_offset_req_1 : boolean;
  signal array_obj_ref_3081_index_offset_ack_1 : boolean;
  signal if_stmt_3216_branch_ack_1 : boolean;
  signal WPIPE_Block3_complete_3336_inst_ack_1 : boolean;
  signal addr_of_3082_final_reg_req_0 : boolean;
  signal addr_of_3082_final_reg_ack_0 : boolean;
  signal type_cast_3240_inst_req_1 : boolean;
  signal if_stmt_3306_branch_req_0 : boolean;
  signal addr_of_3082_final_reg_req_1 : boolean;
  signal ptr_deref_3252_load_0_ack_0 : boolean;
  signal addr_of_3082_final_reg_ack_1 : boolean;
  signal type_cast_2922_inst_ack_1 : boolean;
  signal addr_of_3190_final_reg_ack_1 : boolean;
  signal ptr_deref_3252_load_0_req_0 : boolean;
  signal if_stmt_3216_branch_req_0 : boolean;
  signal ptr_deref_3085_store_0_req_0 : boolean;
  signal ptr_deref_3085_store_0_ack_0 : boolean;
  signal ptr_deref_3085_store_0_req_1 : boolean;
  signal ptr_deref_3085_store_0_ack_1 : boolean;
  signal type_cast_2922_inst_req_1 : boolean;
  signal WPIPE_Block3_complete_3336_inst_req_1 : boolean;
  signal type_cast_3094_inst_req_0 : boolean;
  signal type_cast_3094_inst_ack_0 : boolean;
  signal type_cast_3094_inst_req_1 : boolean;
  signal type_cast_3094_inst_ack_1 : boolean;
  signal phi_stmt_2917_req_0 : boolean;
  signal type_cast_2920_inst_ack_1 : boolean;
  signal type_cast_3282_inst_ack_1 : boolean;
  signal type_cast_3282_inst_req_1 : boolean;
  signal addr_of_3190_final_reg_req_1 : boolean;
  signal type_cast_3158_inst_req_0 : boolean;
  signal type_cast_3158_inst_ack_0 : boolean;
  signal type_cast_3158_inst_req_1 : boolean;
  signal type_cast_3158_inst_ack_1 : boolean;
  signal type_cast_2920_inst_req_1 : boolean;
  signal type_cast_3282_inst_ack_0 : boolean;
  signal type_cast_3282_inst_req_0 : boolean;
  signal type_cast_3201_inst_ack_1 : boolean;
  signal type_cast_3201_inst_req_1 : boolean;
  signal type_cast_3240_inst_ack_0 : boolean;
  signal addr_of_3190_final_reg_ack_0 : boolean;
  signal addr_of_3190_final_reg_req_0 : boolean;
  signal type_cast_3201_inst_ack_0 : boolean;
  signal type_cast_3201_inst_req_0 : boolean;
  signal array_obj_ref_3164_index_offset_req_0 : boolean;
  signal array_obj_ref_3164_index_offset_ack_0 : boolean;
  signal array_obj_ref_3164_index_offset_req_1 : boolean;
  signal array_obj_ref_3164_index_offset_ack_1 : boolean;
  signal WPIPE_Block3_complete_3336_inst_ack_0 : boolean;
  signal WPIPE_Block3_complete_3336_inst_req_0 : boolean;
  signal addr_of_3165_final_reg_req_0 : boolean;
  signal addr_of_3165_final_reg_ack_0 : boolean;
  signal addr_of_3165_final_reg_req_1 : boolean;
  signal addr_of_3165_final_reg_ack_1 : boolean;
  signal ptr_deref_3169_load_0_req_0 : boolean;
  signal ptr_deref_3169_load_0_ack_0 : boolean;
  signal ptr_deref_3169_load_0_req_1 : boolean;
  signal ptr_deref_3169_load_0_ack_1 : boolean;
  signal type_cast_3183_inst_req_0 : boolean;
  signal type_cast_3183_inst_ack_0 : boolean;
  signal type_cast_3183_inst_req_1 : boolean;
  signal type_cast_3183_inst_ack_1 : boolean;
  signal array_obj_ref_3189_index_offset_req_0 : boolean;
  signal array_obj_ref_3189_index_offset_ack_0 : boolean;
  signal array_obj_ref_3189_index_offset_req_1 : boolean;
  signal array_obj_ref_3189_index_offset_ack_1 : boolean;
  signal type_cast_3324_inst_req_0 : boolean;
  signal type_cast_3324_inst_ack_0 : boolean;
  signal type_cast_3324_inst_req_1 : boolean;
  signal type_cast_3324_inst_ack_1 : boolean;
  signal phi_stmt_3319_req_1 : boolean;
  signal type_cast_3316_inst_req_0 : boolean;
  signal type_cast_3316_inst_ack_0 : boolean;
  signal type_cast_3316_inst_req_1 : boolean;
  signal type_cast_3316_inst_ack_1 : boolean;
  signal phi_stmt_3313_req_0 : boolean;
  signal phi_stmt_3325_req_0 : boolean;
  signal type_cast_3322_inst_req_0 : boolean;
  signal type_cast_3322_inst_ack_0 : boolean;
  signal type_cast_3322_inst_req_1 : boolean;
  signal type_cast_3322_inst_ack_1 : boolean;
  signal phi_stmt_3319_req_0 : boolean;
  signal type_cast_3318_inst_req_0 : boolean;
  signal type_cast_3318_inst_ack_0 : boolean;
  signal type_cast_3318_inst_req_1 : boolean;
  signal type_cast_3318_inst_ack_1 : boolean;
  signal phi_stmt_3313_req_1 : boolean;
  signal type_cast_3331_inst_req_0 : boolean;
  signal type_cast_3331_inst_ack_0 : boolean;
  signal type_cast_3331_inst_req_1 : boolean;
  signal type_cast_3331_inst_ack_1 : boolean;
  signal phi_stmt_3325_req_1 : boolean;
  signal phi_stmt_3313_ack_0 : boolean;
  signal phi_stmt_3319_ack_0 : boolean;
  signal phi_stmt_3325_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_D_CP_7327_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_D_CP_7327_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_D_CP_7327_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_D_CP_7327_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_D_CP_7327: Block -- control-path 
    signal zeropad3D_D_CP_7327_elements: BooleanArray(142 downto 0);
    -- 
  begin -- 
    zeropad3D_D_CP_7327_elements(0) <= zeropad3D_D_CP_7327_start;
    zeropad3D_D_CP_7327_symbol <= zeropad3D_D_CP_7327_elements(94);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2717/$entry
      -- CP-element group 0: 	 branch_block_stmt_2717/branch_block_stmt_2717__entry__
      -- CP-element group 0: 	 branch_block_stmt_2717/assign_stmt_2720__entry__
      -- CP-element group 0: 	 branch_block_stmt_2717/assign_stmt_2720/$entry
      -- CP-element group 0: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Sample/rr
      -- 
    rr_7405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(0), ack => RPIPE_Block3_starting_2719_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	142 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	104 
    -- CP-element group 1: 	106 
    -- CP-element group 1: 	107 
    -- CP-element group 1: 	109 
    -- CP-element group 1: 	110 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/merge_stmt_3312__exit__
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/$entry
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/$entry
      -- 
    rr_8652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(1), ack => type_cast_2928_inst_req_0); -- 
    rr_8629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(1), ack => type_cast_2922_inst_req_0); -- 
    cr_8657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(1), ack => type_cast_2928_inst_req_1); -- 
    cr_8680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(1), ack => type_cast_2935_inst_req_1); -- 
    rr_8675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(1), ack => type_cast_2935_inst_req_0); -- 
    cr_8634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(1), ack => type_cast_2922_inst_req_1); -- 
    zeropad3D_D_CP_7327_elements(1) <= zeropad3D_D_CP_7327_elements(142);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Update/cr
      -- 
    ra_7406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2719_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(2)); -- 
    cr_7410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(2), ack => RPIPE_Block3_starting_2719_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	18 
    -- CP-element group 3: 	19 
    -- CP-element group 3: 	14 
    -- CP-element group 3: 	9 
    -- CP-element group 3: 	11 
    -- CP-element group 3: 	13 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	15 
    -- CP-element group 3: 	16 
    -- CP-element group 3: 	17 
    -- CP-element group 3: 	21 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	7 
    -- CP-element group 3:  members (158) 
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2720__exit__
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914__entry__
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2720/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2720/RPIPE_Block3_starting_2719_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Update/cr
      -- 
    ca_7411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2719_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(3)); -- 
    cr_7541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => type_cast_2764_inst_req_1); -- 
    cr_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2754_load_0_req_1); -- 
    rr_7511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2754_load_0_req_0); -- 
    cr_7458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2732_load_0_req_1); -- 
    rr_7558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => LOAD_pad_2767_load_0_req_0); -- 
    cr_7569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => LOAD_pad_2767_load_0_req_1); -- 
    cr_7477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => type_cast_2742_inst_req_1); -- 
    rr_7608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2779_load_0_req_0); -- 
    rr_7447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2732_load_0_req_0); -- 
    cr_7619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2779_load_0_req_1); -- 
    rr_7658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2791_load_0_req_0); -- 
    cr_7669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2791_load_0_req_1); -- 
    rr_7708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2803_load_0_req_0); -- 
    cr_7719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => ptr_deref_2803_load_0_req_1); -- 
    cr_7738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(3), ack => type_cast_2857_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/word_access_start/word_0/ra
      -- CP-element group 4: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Sample/word_access_start/$exit
      -- 
    ra_7448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (12) 
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/word_access_complete/word_0/ca
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/ptr_deref_2732_Merge/merge_req
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/ptr_deref_2732_Merge/$entry
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/ptr_deref_2732_Merge/$exit
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_Update/ptr_deref_2732_Merge/merge_ack
      -- CP-element group 5: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2732_update_completed_
      -- 
    ca_7459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(5)); -- 
    rr_7472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(5), ack => type_cast_2742_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Sample/ra
      -- 
    ra_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2742_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	3 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	22 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2742_Update/$exit
      -- 
    ca_7478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2742_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Sample/word_access_start/word_0/$exit
      -- 
    ra_7512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2754_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	3 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (12) 
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/ptr_deref_2754_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/ptr_deref_2754_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/ptr_deref_2754_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/ptr_deref_2754_Merge/merge_ack
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2754_Update/$exit
      -- 
    ca_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2754_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(9)); -- 
    rr_7536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(9), ack => type_cast_2764_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Sample/ra
      -- 
    ra_7537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2764_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	22 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2764_Update/ca
      -- 
    ca_7542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2764_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/word_access_start/word_0/ra
      -- CP-element group 12: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Sample/word_access_start/$exit
      -- 
    ra_7559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2767_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	20 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/LOAD_pad_2767_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/LOAD_pad_2767_Merge/merge_ack
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/LOAD_pad_2767_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/LOAD_pad_2767_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/LOAD_pad_2767_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Sample/rr
      -- 
    ca_7570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2767_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(13)); -- 
    rr_7733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(13), ack => type_cast_2857_inst_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	3 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Sample/word_access_start/word_0/ra
      -- 
    ra_7609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2779_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/ptr_deref_2779_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/ptr_deref_2779_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/ptr_deref_2779_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2779_Update/ptr_deref_2779_Merge/merge_ack
      -- 
    ca_7620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2779_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Sample/word_access_start/word_0/ra
      -- 
    ra_7659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2791_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	22 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/ptr_deref_2791_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/ptr_deref_2791_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/ptr_deref_2791_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2791_Update/ptr_deref_2791_Merge/merge_ack
      -- 
    ca_7670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2791_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	3 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/word_access_start/$exit
      -- CP-element group 18: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Sample/word_access_start/word_0/ra
      -- 
    ra_7709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2803_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	3 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/word_access_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/ptr_deref_2803_Merge/$entry
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/ptr_deref_2803_Merge/$exit
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/ptr_deref_2803_Merge/merge_req
      -- CP-element group 19: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/ptr_deref_2803_Update/ptr_deref_2803_Merge/merge_ack
      -- 
    ca_7720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2803_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	13 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Sample/ra
      -- 
    ra_7734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	3 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/type_cast_2857_Update/ca
      -- 
    ca_7739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(21)); -- 
    -- CP-element group 22:  join  fork  transition  place  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	11 
    -- CP-element group 22: 	15 
    -- CP-element group 22: 	17 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	95 
    -- CP-element group 22: 	96 
    -- CP-element group 22: 	98 
    -- CP-element group 22: 	99 
    -- CP-element group 22: 	101 
    -- CP-element group 22:  members (22) 
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Update/cr
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2929/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914__exit__
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody
      -- CP-element group 22: 	 branch_block_stmt_2717/assign_stmt_2729_to_assign_stmt_2914/$exit
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/$entry
      -- CP-element group 22: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Update/cr
      -- 
    cr_8600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(22), ack => type_cast_2926_inst_req_1); -- 
    rr_8572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(22), ack => type_cast_2920_inst_req_0); -- 
    rr_8595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(22), ack => type_cast_2926_inst_req_0); -- 
    cr_8577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(22), ack => type_cast_2920_inst_req_1); -- 
    zeropad3D_D_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(19) & zeropad3D_D_CP_7327_elements(11) & zeropad3D_D_CP_7327_elements(15) & zeropad3D_D_CP_7327_elements(17) & zeropad3D_D_CP_7327_elements(21) & zeropad3D_D_CP_7327_elements(7);
      gj_zeropad3D_D_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	117 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Sample/ra
      -- 
    ra_7751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2940_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(23)); -- 
    -- CP-element group 24:  branch  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	117 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (13) 
      -- CP-element group 24: 	 branch_block_stmt_2717/R_cmp_2950_place
      -- CP-element group 24: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948__exit__
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949__entry__
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949_dead_link/$entry
      -- CP-element group 24: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/$exit
      -- CP-element group 24: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949_eval_test/$entry
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949_eval_test/$exit
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949_eval_test/branch_req
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949_if_link/$entry
      -- CP-element group 24: 	 branch_block_stmt_2717/if_stmt_2949_else_link/$entry
      -- 
    ca_7756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2940_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(24)); -- 
    branch_req_7764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(24), ack => if_stmt_2949_branch_req_0); -- 
    -- CP-element group 25:  transition  place  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	118 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2717/whilex_xbody_ifx_xthen
      -- CP-element group 25: 	 branch_block_stmt_2717/if_stmt_2949_if_link/$exit
      -- CP-element group 25: 	 branch_block_stmt_2717/if_stmt_2949_if_link/if_choice_transition
      -- CP-element group 25: 	 branch_block_stmt_2717/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 25: 	 branch_block_stmt_2717/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_7769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2949_branch_ack_1, ack => zeropad3D_D_CP_7327_elements(25)); -- 
    -- CP-element group 26:  merge  transition  place  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (11) 
      -- CP-element group 26: 	 branch_block_stmt_2717/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 26: 	 branch_block_stmt_2717/merge_stmt_2955_PhiReqMerge
      -- CP-element group 26: 	 branch_block_stmt_2717/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- CP-element group 26: 	 branch_block_stmt_2717/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 26: 	 branch_block_stmt_2717/merge_stmt_2955_PhiAck/$entry
      -- CP-element group 26: 	 branch_block_stmt_2717/merge_stmt_2955_PhiAck/$exit
      -- CP-element group 26: 	 branch_block_stmt_2717/merge_stmt_2955_PhiAck/dummy
      -- CP-element group 26: 	 branch_block_stmt_2717/merge_stmt_2955__exit__
      -- CP-element group 26: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977__entry__
      -- CP-element group 26: 	 branch_block_stmt_2717/if_stmt_2949_else_link/$exit
      -- CP-element group 26: 	 branch_block_stmt_2717/if_stmt_2949_else_link/else_choice_transition
      -- 
    else_choice_transition_7773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2949_branch_ack_0, ack => zeropad3D_D_CP_7327_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (27) 
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_update_start_
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_address_calculated
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_word_address_calculated
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_root_address_calculated
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_address_resized
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_addr_resize/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_addr_resize/$exit
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_addr_resize/base_resize_req
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_addr_resize/base_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_plus_offset/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_plus_offset/$exit
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_plus_offset/sum_rename_req
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_base_plus_offset/sum_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_word_addrgen/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_word_addrgen/$exit
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_word_addrgen/root_register_req
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_word_addrgen/root_register_ack
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/word_access_start/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/word_access_start/word_0/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/word_access_start/word_0/rr
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/word_access_complete/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/word_access_complete/word_0/$entry
      -- CP-element group 27: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/word_access_complete/word_0/cr
      -- 
    cr_7822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(27), ack => ptr_deref_2966_load_0_req_1); -- 
    rr_7811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(27), ack => ptr_deref_2966_load_0_req_0); -- 
    zeropad3D_D_CP_7327_elements(27) <= zeropad3D_D_CP_7327_elements(26);
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/word_access_start/$exit
      -- CP-element group 28: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/word_access_start/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Sample/word_access_start/word_0/ra
      -- 
    ra_7812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2966_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(28)); -- 
    -- CP-element group 29:  branch  transition  place  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (19) 
      -- CP-element group 29: 	 branch_block_stmt_2717/R_cmp52_2979_place
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977__exit__
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978__entry__
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/$exit
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/word_access_complete/$exit
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/word_access_complete/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/word_access_complete/word_0/ca
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/ptr_deref_2966_Merge/$entry
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/ptr_deref_2966_Merge/$exit
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/ptr_deref_2966_Merge/merge_req
      -- CP-element group 29: 	 branch_block_stmt_2717/assign_stmt_2963_to_assign_stmt_2977/ptr_deref_2966_Update/ptr_deref_2966_Merge/merge_ack
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978_dead_link/$entry
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978_eval_test/$entry
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978_eval_test/$exit
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978_eval_test/branch_req
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978_if_link/$entry
      -- CP-element group 29: 	 branch_block_stmt_2717/if_stmt_2978_else_link/$entry
      -- 
    ca_7823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2966_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(29)); -- 
    branch_req_7836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(29), ack => if_stmt_2978_branch_req_0); -- 
    -- CP-element group 30:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (18) 
      -- CP-element group 30: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse54
      -- CP-element group 30: 	 branch_block_stmt_2717/merge_stmt_2984_PhiReqMerge
      -- CP-element group 30: 	 branch_block_stmt_2717/merge_stmt_2984__exit__
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996__entry__
      -- CP-element group 30: 	 branch_block_stmt_2717/if_stmt_2978_if_link/$exit
      -- CP-element group 30: 	 branch_block_stmt_2717/if_stmt_2978_if_link/if_choice_transition
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/$entry
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse54_PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse54_PhiReq/$exit
      -- CP-element group 30: 	 branch_block_stmt_2717/merge_stmt_2984_PhiAck/$entry
      -- CP-element group 30: 	 branch_block_stmt_2717/merge_stmt_2984_PhiAck/$exit
      -- CP-element group 30: 	 branch_block_stmt_2717/merge_stmt_2984_PhiAck/dummy
      -- 
    if_choice_transition_7841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2978_branch_ack_1, ack => zeropad3D_D_CP_7327_elements(30)); -- 
    rr_7858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(30), ack => type_cast_2988_inst_req_0); -- 
    cr_7863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(30), ack => type_cast_2988_inst_req_1); -- 
    -- CP-element group 31:  transition  place  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	118 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 31: 	 branch_block_stmt_2717/if_stmt_2978_else_link/$exit
      -- CP-element group 31: 	 branch_block_stmt_2717/if_stmt_2978_else_link/else_choice_transition
      -- CP-element group 31: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_7845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2978_branch_ack_0, ack => zeropad3D_D_CP_7327_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Sample/ra
      -- 
    ra_7859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2988_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(32)); -- 
    -- CP-element group 33:  branch  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (13) 
      -- CP-element group 33: 	 branch_block_stmt_2717/R_cmp59_2998_place
      -- CP-element group 33: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996__exit__
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997__entry__
      -- CP-element group 33: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/$exit
      -- CP-element group 33: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2717/assign_stmt_2989_to_assign_stmt_2996/type_cast_2988_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997_dead_link/$entry
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997_eval_test/$entry
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997_eval_test/$exit
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997_eval_test/branch_req
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997_if_link/$entry
      -- CP-element group 33: 	 branch_block_stmt_2717/if_stmt_2997_else_link/$entry
      -- 
    ca_7864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2988_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(33)); -- 
    branch_req_7872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(33), ack => if_stmt_2997_branch_req_0); -- 
    -- CP-element group 34:  transition  place  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	118 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse54_ifx_xthen
      -- CP-element group 34: 	 branch_block_stmt_2717/if_stmt_2997_if_link/$exit
      -- CP-element group 34: 	 branch_block_stmt_2717/if_stmt_2997_if_link/if_choice_transition
      -- CP-element group 34: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_7877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2997_branch_ack_1, ack => zeropad3D_D_CP_7327_elements(34)); -- 
    -- CP-element group 35:  merge  transition  place  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (11) 
      -- CP-element group 35: 	 branch_block_stmt_2717/merge_stmt_3003_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_2717/merge_stmt_3003__exit__
      -- CP-element group 35: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025__entry__
      -- CP-element group 35: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse54_lorx_xlhsx_xfalse61_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_2717/if_stmt_2997_else_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_2717/if_stmt_2997_else_link/else_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse54_lorx_xlhsx_xfalse61
      -- CP-element group 35: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse54_lorx_xlhsx_xfalse61_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_2717/merge_stmt_3003_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_2717/merge_stmt_3003_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_2717/merge_stmt_3003_PhiAck/dummy
      -- 
    else_choice_transition_7881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2997_branch_ack_0, ack => zeropad3D_D_CP_7327_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (27) 
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_update_start_
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_address_calculated
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_word_address_calculated
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_root_address_calculated
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_address_resized
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_addr_resize/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_addr_resize/$exit
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_addr_resize/base_resize_req
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_addr_resize/base_resize_ack
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_plus_offset/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_plus_offset/$exit
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_plus_offset/sum_rename_req
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_base_plus_offset/sum_rename_ack
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_word_addrgen/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_word_addrgen/$exit
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_word_addrgen/root_register_req
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_word_addrgen/root_register_ack
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/word_access_start/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/word_access_start/word_0/rr
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/word_access_complete/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/word_access_complete/word_0/$entry
      -- CP-element group 36: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/word_access_complete/word_0/cr
      -- 
    cr_7930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(36), ack => ptr_deref_3014_load_0_req_1); -- 
    rr_7919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(36), ack => ptr_deref_3014_load_0_req_0); -- 
    zeropad3D_D_CP_7327_elements(36) <= zeropad3D_D_CP_7327_elements(35);
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/word_access_start/$exit
      -- CP-element group 37: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Sample/word_access_start/word_0/ra
      -- 
    ra_7920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3014_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (19) 
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025__exit__
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026__entry__
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/$exit
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/word_access_complete/$exit
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/word_access_complete/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/word_access_complete/word_0/ca
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/ptr_deref_3014_Merge/$entry
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/ptr_deref_3014_Merge/$exit
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/ptr_deref_3014_Merge/merge_req
      -- CP-element group 38: 	 branch_block_stmt_2717/assign_stmt_3011_to_assign_stmt_3025/ptr_deref_3014_Update/ptr_deref_3014_Merge/merge_ack
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026_eval_test/branch_req
      -- CP-element group 38: 	 branch_block_stmt_2717/R_cmp68_3027_place
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026_if_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_2717/if_stmt_3026_else_link/$entry
      -- 
    ca_7931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3014_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(38)); -- 
    branch_req_7944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(38), ack => if_stmt_3026_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_2717/merge_stmt_3090_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/merge_stmt_3090__exit__
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195__entry__
      -- CP-element group 39: 	 branch_block_stmt_2717/if_stmt_3026_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_2717/if_stmt_3026_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse61_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_complete/req
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_complete/req
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse61_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse61_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_2717/merge_stmt_3090_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_2717/merge_stmt_3090_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_2717/merge_stmt_3090_PhiAck/dummy
      -- 
    if_choice_transition_7949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3026_branch_ack_1, ack => zeropad3D_D_CP_7327_elements(39)); -- 
    cr_8332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => ptr_deref_3193_store_0_req_1); -- 
    rr_8107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => type_cast_3094_inst_req_0); -- 
    cr_8112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => type_cast_3094_inst_req_1); -- 
    req_8282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => addr_of_3190_final_reg_req_1); -- 
    cr_8126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => type_cast_3158_inst_req_1); -- 
    req_8157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => array_obj_ref_3164_index_offset_req_1); -- 
    req_8172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => addr_of_3165_final_reg_req_1); -- 
    cr_8217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => ptr_deref_3169_load_0_req_1); -- 
    cr_8236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => type_cast_3183_inst_req_1); -- 
    req_8267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(39), ack => array_obj_ref_3189_index_offset_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	118 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_2717/if_stmt_3026_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_2717/if_stmt_3026_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse61_ifx_xthen
      -- CP-element group 40: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse61_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_2717/lorx_xlhsx_xfalse61_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_7953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3026_branch_ack_0, ack => zeropad3D_D_CP_7327_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	118 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Sample/ra
      -- 
    ra_7967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3036_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	118 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Update/ca
      -- 
    ca_7972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3036_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	118 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Sample/ra
      -- 
    ra_7981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3041_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	118 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Update/ca
      -- 
    ca_7986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3041_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Sample/rr
      -- 
    rr_7994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(45), ack => type_cast_3075_inst_req_0); -- 
    zeropad3D_D_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(42) & zeropad3D_D_CP_7327_elements(44);
      gj_zeropad3D_D_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Sample/ra
      -- 
    ra_7995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3075_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	118 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_computed_1
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Sample/req
      -- 
    ca_8000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3075_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(47)); -- 
    req_8025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(47), ack => array_obj_ref_3081_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Sample/ack
      -- 
    ack_8026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3081_index_offset_ack_0, ack => zeropad3D_D_CP_7327_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	118 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_request/req
      -- 
    ack_8031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3081_index_offset_ack_1, ack => zeropad3D_D_CP_7327_elements(49)); -- 
    req_8040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(49), ack => addr_of_3082_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_request/$exit
      -- CP-element group 50: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_request/ack
      -- 
    ack_8041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3082_final_reg_ack_0, ack => zeropad3D_D_CP_7327_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	118 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_word_addrgen/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/ptr_deref_3085_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/ptr_deref_3085_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/ptr_deref_3085_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/ptr_deref_3085_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/word_access_start/word_0/rr
      -- 
    ack_8046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3082_final_reg_ack_1, ack => zeropad3D_D_CP_7327_elements(51)); -- 
    rr_8084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(51), ack => ptr_deref_3085_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Sample/word_access_start/word_0/ra
      -- 
    ra_8085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3085_store_0_ack_0, ack => zeropad3D_D_CP_7327_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	118 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/word_access_complete/word_0/ca
      -- 
    ca_8096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3085_store_0_ack_1, ack => zeropad3D_D_CP_7327_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	48 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	119 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088__exit__
      -- CP-element group 54: 	 branch_block_stmt_2717/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/$exit
      -- CP-element group 54: 	 branch_block_stmt_2717/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2717/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(48) & zeropad3D_D_CP_7327_elements(53);
      gj_zeropad3D_D_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Sample/ra
      -- 
    ra_8108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3094_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3094_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Sample/rr
      -- 
    ca_8113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3094_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(56)); -- 
    rr_8121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(56), ack => type_cast_3158_inst_req_0); -- 
    rr_8231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(56), ack => type_cast_3183_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Sample/ra
      -- 
    ra_8122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3158_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3158_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Sample/req
      -- 
    ca_8127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3158_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(58)); -- 
    req_8152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(58), ack => array_obj_ref_3164_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Sample/ack
      -- 
    ack_8153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3164_index_offset_ack_0, ack => zeropad3D_D_CP_7327_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3164_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_request/req
      -- 
    ack_8158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3164_index_offset_ack_1, ack => zeropad3D_D_CP_7327_elements(60)); -- 
    req_8167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(60), ack => addr_of_3165_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_request/ack
      -- 
    ack_8168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3165_final_reg_ack_0, ack => zeropad3D_D_CP_7327_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3165_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/word_access_start/word_0/rr
      -- 
    ack_8173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3165_final_reg_ack_1, ack => zeropad3D_D_CP_7327_elements(62)); -- 
    rr_8206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(62), ack => ptr_deref_3169_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Sample/word_access_start/word_0/ra
      -- 
    ra_8207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3169_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/ptr_deref_3169_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/ptr_deref_3169_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/ptr_deref_3169_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3169_Update/ptr_deref_3169_Merge/merge_ack
      -- 
    ca_8218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3169_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Sample/ra
      -- 
    ra_8232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3183_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/type_cast_3183_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_computed_1
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Sample/req
      -- 
    ca_8237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3183_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(66)); -- 
    req_8262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(66), ack => array_obj_ref_3189_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Sample/ack
      -- 
    ack_8263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3189_index_offset_ack_0, ack => zeropad3D_D_CP_7327_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_request/req
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/array_obj_ref_3189_base_plus_offset/sum_rename_ack
      -- 
    ack_8268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3189_index_offset_ack_1, ack => zeropad3D_D_CP_7327_elements(68)); -- 
    req_8277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(68), ack => addr_of_3190_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_request/ack
      -- CP-element group 69: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_sample_completed_
      -- 
    ack_8278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3190_final_reg_ack_0, ack => zeropad3D_D_CP_7327_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_word_addrgen/root_register_ack
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/addr_of_3190_update_completed_
      -- 
    ack_8283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3190_final_reg_ack_1, ack => zeropad3D_D_CP_7327_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/word_access_start/word_0/rr
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/ptr_deref_3193_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/ptr_deref_3193_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/ptr_deref_3193_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/ptr_deref_3193_Split/$entry
      -- 
    rr_8321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(71), ack => ptr_deref_3193_store_0_req_0); -- 
    zeropad3D_D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(64) & zeropad3D_D_CP_7327_elements(70);
      gj_zeropad3D_D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/word_access_start/word_0/ra
      -- CP-element group 72: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Sample/word_access_start/$exit
      -- 
    ra_8322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3193_store_0_ack_0, ack => zeropad3D_D_CP_7327_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/word_access_complete/word_0/ca
      -- CP-element group 73: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/ptr_deref_3193_Update/$exit
      -- 
    ca_8333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3193_store_0_ack_1, ack => zeropad3D_D_CP_7327_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	119 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195__exit__
      -- CP-element group 74: 	 branch_block_stmt_2717/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_2717/assign_stmt_3095_to_assign_stmt_3195/$exit
      -- CP-element group 74: 	 branch_block_stmt_2717/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2717/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(59) & zeropad3D_D_CP_7327_elements(67) & zeropad3D_D_CP_7327_elements(73);
      gj_zeropad3D_D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	119 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_sample_completed_
      -- 
    ra_8345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3201_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	119 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215__exit__
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216__entry__
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216_else_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_2717/R_cmp137_3217_place
      -- CP-element group 76: 	 branch_block_stmt_2717/if_stmt_3216_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/$exit
      -- 
    ca_8350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3201_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(76)); -- 
    branch_req_8358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(76), ack => if_stmt_3216_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	128 
    -- CP-element group 77: 	129 
    -- CP-element group 77: 	131 
    -- CP-element group 77: 	132 
    -- CP-element group 77: 	134 
    -- CP-element group 77: 	135 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_2717/merge_stmt_3222__exit__
      -- CP-element group 77: 	 branch_block_stmt_2717/assign_stmt_3228__entry__
      -- CP-element group 77: 	 branch_block_stmt_2717/assign_stmt_3228__exit__
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xend_ifx_xthen139
      -- CP-element group 77: 	 branch_block_stmt_2717/assign_stmt_3228/$exit
      -- CP-element group 77: 	 branch_block_stmt_2717/assign_stmt_3228/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/if_stmt_3216_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_2717/if_stmt_3216_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xend_ifx_xthen139_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xend_ifx_xthen139_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_2717/merge_stmt_3222_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_2717/merge_stmt_3222_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/merge_stmt_3222_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_2717/merge_stmt_3222_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3216_branch_ack_1, ack => zeropad3D_D_CP_7327_elements(77)); -- 
    rr_8865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(77), ack => type_cast_3322_inst_req_0); -- 
    cr_8870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(77), ack => type_cast_3322_inst_req_1); -- 
    rr_8888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(77), ack => type_cast_3318_inst_req_0); -- 
    cr_8893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(77), ack => type_cast_3318_inst_req_1); -- 
    rr_8911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(77), ack => type_cast_3331_inst_req_0); -- 
    cr_8916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(77), ack => type_cast_3331_inst_req_1); -- 
    -- CP-element group 78:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	81 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	85 
    -- CP-element group 78: 	87 
    -- CP-element group 78: 	88 
    -- CP-element group 78: 	89 
    -- CP-element group 78:  members (76) 
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/word_access_complete/word_0/cr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/word_access_start/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/word_access_start/word_0/rr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_word_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_root_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_address_resized
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_addr_resize/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_addr_resize/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_addr_resize/base_resize_req
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_addr_resize/base_resize_ack
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/word_access_complete/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/merge_stmt_3230__exit__
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305__entry__
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_word_addrgen/root_register_ack
      -- CP-element group 78: 	 branch_block_stmt_2717/ifx_xend_ifx_xelse144
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_word_addrgen/root_register_req
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_word_addrgen/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_word_addrgen/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_plus_offset/sum_rename_ack
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_plus_offset/sum_rename_req
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_plus_offset/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/word_access_complete/word_0/cr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_plus_offset/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_addr_resize/base_resize_ack
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_addr_resize/base_resize_req
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_addr_resize/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_addr_resize/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_address_resized
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_root_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/if_stmt_3216_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_2717/if_stmt_3216_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/word_access_complete/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/word_access_complete/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_word_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_base_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/word_access_start/word_0/rr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/word_access_start/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/word_access_start/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/word_access_complete/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/word_access_start/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_word_addrgen/root_register_ack
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_word_addrgen/root_register_req
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_word_addrgen/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_word_addrgen/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_plus_offset/sum_rename_ack
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_plus_offset/sum_rename_req
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_plus_offset/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_base_plus_offset/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/ifx_xend_ifx_xelse144_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/ifx_xend_ifx_xelse144_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/merge_stmt_3230_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2717/merge_stmt_3230_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2717/merge_stmt_3230_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2717/merge_stmt_3230_PhiAck/dummy
      -- 
    else_choice_transition_8367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3216_branch_ack_0, ack => zeropad3D_D_CP_7327_elements(78)); -- 
    cr_8511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => ptr_deref_3294_load_0_req_1); -- 
    rr_8500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => ptr_deref_3294_load_0_req_0); -- 
    cr_8452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => type_cast_3266_inst_req_1); -- 
    rr_8383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => type_cast_3240_inst_req_0); -- 
    cr_8433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => ptr_deref_3252_load_0_req_1); -- 
    cr_8388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => type_cast_3240_inst_req_1); -- 
    rr_8422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => ptr_deref_3252_load_0_req_0); -- 
    cr_8466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(78), ack => type_cast_3282_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Sample/ra
      -- 
    ra_8384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3240_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3240_Update/$exit
      -- 
    ca_8389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3240_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/word_access_start/word_0/ra
      -- CP-element group 81: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/word_access_start/$exit
      -- CP-element group 81: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Sample/$exit
      -- 
    ra_8423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3252_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/ptr_deref_3252_Merge/merge_ack
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/ptr_deref_3252_Merge/merge_req
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/ptr_deref_3252_Merge/$exit
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/ptr_deref_3252_Merge/$entry
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/word_access_complete/word_0/ca
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/word_access_complete/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/word_access_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3252_Update/$exit
      -- 
    ca_8434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3252_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_sample_start_
      -- 
    rr_8447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(83), ack => type_cast_3266_inst_req_0); -- 
    zeropad3D_D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(80) & zeropad3D_D_CP_7327_elements(82);
      gj_zeropad3D_D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_sample_completed_
      -- 
    ra_8448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3266_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	78 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3266_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Sample/$entry
      -- 
    ca_8453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3266_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(85)); -- 
    rr_8461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(85), ack => type_cast_3282_inst_req_0); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Sample/$exit
      -- 
    ra_8462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3282_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	78 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/type_cast_3282_update_completed_
      -- 
    ca_8467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3282_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	78 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/word_access_start/word_0/ra
      -- CP-element group 88: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_sample_completed_
      -- 
    ra_8501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_load_0_ack_0, ack => zeropad3D_D_CP_7327_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	78 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (9) 
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/word_access_complete/word_0/ca
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/ptr_deref_3294_Merge/$entry
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/word_access_complete/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/ptr_deref_3294_Merge/merge_ack
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/ptr_deref_3294_Merge/merge_req
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/ptr_deref_3294_Update/ptr_deref_3294_Merge/$exit
      -- 
    ca_8512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_load_0_ack_1, ack => zeropad3D_D_CP_7327_elements(89)); -- 
    -- CP-element group 90:  branch  join  transition  place  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (10) 
      -- CP-element group 90: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305__exit__
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306__entry__
      -- CP-element group 90: 	 branch_block_stmt_2717/R_cmp166_3307_place
      -- CP-element group 90: 	 branch_block_stmt_2717/assign_stmt_3236_to_assign_stmt_3305/$exit
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306_else_link/$entry
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306_if_link/$entry
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306_eval_test/branch_req
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306_eval_test/$exit
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306_eval_test/$entry
      -- CP-element group 90: 	 branch_block_stmt_2717/if_stmt_3306_dead_link/$entry
      -- 
    branch_req_8525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(90), ack => if_stmt_3306_branch_req_0); -- 
    zeropad3D_D_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(87) & zeropad3D_D_CP_7327_elements(89);
      gj_zeropad3D_D_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  place  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (15) 
      -- CP-element group 91: 	 branch_block_stmt_2717/ifx_xelse144_whilex_xend
      -- CP-element group 91: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2717/merge_stmt_3334__exit__
      -- CP-element group 91: 	 branch_block_stmt_2717/assign_stmt_3338__entry__
      -- CP-element group 91: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2717/assign_stmt_3338/$entry
      -- CP-element group 91: 	 branch_block_stmt_2717/if_stmt_3306_if_link/if_choice_transition
      -- CP-element group 91: 	 branch_block_stmt_2717/if_stmt_3306_if_link/$exit
      -- CP-element group 91: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Sample/req
      -- CP-element group 91: 	 branch_block_stmt_2717/ifx_xelse144_whilex_xend_PhiReq/$entry
      -- CP-element group 91: 	 branch_block_stmt_2717/ifx_xelse144_whilex_xend_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_2717/merge_stmt_3334_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_2717/merge_stmt_3334_PhiAck/$entry
      -- CP-element group 91: 	 branch_block_stmt_2717/merge_stmt_3334_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_2717/merge_stmt_3334_PhiAck/dummy
      -- 
    if_choice_transition_8530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3306_branch_ack_1, ack => zeropad3D_D_CP_7327_elements(91)); -- 
    req_8547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(91), ack => WPIPE_Block3_complete_3336_inst_req_0); -- 
    -- CP-element group 92:  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	120 
    -- CP-element group 92: 	121 
    -- CP-element group 92: 	123 
    -- CP-element group 92: 	124 
    -- CP-element group 92: 	126 
    -- CP-element group 92:  members (22) 
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174
      -- CP-element group 92: 	 branch_block_stmt_2717/if_stmt_3306_else_link/else_choice_transition
      -- CP-element group 92: 	 branch_block_stmt_2717/if_stmt_3306_else_link/$exit
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3325/$entry
      -- CP-element group 92: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/$entry
      -- 
    else_choice_transition_8534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3306_branch_ack_0, ack => zeropad3D_D_CP_7327_elements(92)); -- 
    rr_8808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(92), ack => type_cast_3324_inst_req_0); -- 
    cr_8813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(92), ack => type_cast_3324_inst_req_1); -- 
    rr_8831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(92), ack => type_cast_3316_inst_req_0); -- 
    cr_8836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(92), ack => type_cast_3316_inst_req_1); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_update_start_
      -- CP-element group 93: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Update/req
      -- CP-element group 93: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Sample/ack
      -- 
    ack_8548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_complete_3336_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(93)); -- 
    req_8552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(93), ack => WPIPE_Block3_complete_3336_inst_req_1); -- 
    -- CP-element group 94:  transition  place  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (16) 
      -- CP-element group 94: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_update_completed_
      -- CP-element group 94: 	 $exit
      -- CP-element group 94: 	 branch_block_stmt_2717/$exit
      -- CP-element group 94: 	 branch_block_stmt_2717/branch_block_stmt_2717__exit__
      -- CP-element group 94: 	 branch_block_stmt_2717/assign_stmt_3338__exit__
      -- CP-element group 94: 	 branch_block_stmt_2717/return__
      -- CP-element group 94: 	 branch_block_stmt_2717/merge_stmt_3340__exit__
      -- CP-element group 94: 	 branch_block_stmt_2717/assign_stmt_3338/$exit
      -- CP-element group 94: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_2717/assign_stmt_3338/WPIPE_Block3_complete_3336_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2717/return___PhiReq/$entry
      -- CP-element group 94: 	 branch_block_stmt_2717/return___PhiReq/$exit
      -- CP-element group 94: 	 branch_block_stmt_2717/merge_stmt_3340_PhiReqMerge
      -- CP-element group 94: 	 branch_block_stmt_2717/merge_stmt_3340_PhiAck/$entry
      -- CP-element group 94: 	 branch_block_stmt_2717/merge_stmt_3340_PhiAck/$exit
      -- CP-element group 94: 	 branch_block_stmt_2717/merge_stmt_3340_PhiAck/dummy
      -- 
    ack_8553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_complete_3336_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	22 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Sample/ra
      -- 
    ra_8573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2920_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	22 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Update/ca
      -- CP-element group 96: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/Update/$exit
      -- 
    ca_8578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2920_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	102 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/$exit
      -- CP-element group 97: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2920/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/$exit
      -- CP-element group 97: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_req
      -- 
    phi_stmt_2917_req_8579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2917_req_8579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(97), ack => phi_stmt_2917_req_0); -- 
    zeropad3D_D_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(95) & zeropad3D_D_CP_7327_elements(96);
      gj_zeropad3D_D_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	22 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Sample/$exit
      -- 
    ra_8596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2926_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	22 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Update/ca
      -- CP-element group 99: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/Update/$exit
      -- 
    ca_8601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2926_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_req
      -- CP-element group 100: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2926/$exit
      -- CP-element group 100: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2923/$exit
      -- 
    phi_stmt_2923_req_8602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2923_req_8602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(100), ack => phi_stmt_2923_req_0); -- 
    zeropad3D_D_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(98) & zeropad3D_D_CP_7327_elements(99);
      gj_zeropad3D_D_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	22 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_req
      -- CP-element group 101: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2933_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2929/$exit
      -- CP-element group 101: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/$exit
      -- 
    phi_stmt_2929_req_8610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2929_req_8610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(101), ack => phi_stmt_2929_req_0); -- 
    -- Element group zeropad3D_D_CP_7327_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => zeropad3D_D_CP_7327_elements(22), ack => zeropad3D_D_CP_7327_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	97 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	113 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2717/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(97) & zeropad3D_D_CP_7327_elements(100) & zeropad3D_D_CP_7327_elements(101);
      gj_zeropad3D_D_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Sample/$exit
      -- 
    ra_8630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2922_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	1 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/Update/$exit
      -- 
    ca_8635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2922_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/$exit
      -- CP-element group 105: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/$exit
      -- CP-element group 105: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/type_cast_2922/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2917/phi_stmt_2917_req
      -- 
    phi_stmt_2917_req_8636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2917_req_8636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(105), ack => phi_stmt_2917_req_1); -- 
    zeropad3D_D_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(103) & zeropad3D_D_CP_7327_elements(104);
      gj_zeropad3D_D_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Sample/$exit
      -- 
    ra_8653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2928_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	1 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Update/ca
      -- CP-element group 107: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/Update/$exit
      -- 
    ca_8658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2928_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_req
      -- CP-element group 108: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/phi_stmt_2923_sources/type_cast_2928/$exit
      -- CP-element group 108: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2923/$exit
      -- 
    phi_stmt_2923_req_8659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2923_req_8659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(108), ack => phi_stmt_2923_req_1); -- 
    zeropad3D_D_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(106) & zeropad3D_D_CP_7327_elements(107);
      gj_zeropad3D_D_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	1 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Sample/ra
      -- 
    ra_8676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2935_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	1 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/Update/ca
      -- 
    ca_8681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2935_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_req
      -- CP-element group 111: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/$exit
      -- CP-element group 111: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/$exit
      -- CP-element group 111: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_2929/phi_stmt_2929_sources/type_cast_2935/SplitProtocol/$exit
      -- 
    phi_stmt_2929_req_8682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2929_req_8682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(111), ack => phi_stmt_2929_req_1); -- 
    zeropad3D_D_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(109) & zeropad3D_D_CP_7327_elements(110);
      gj_zeropad3D_D_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2717/ifx_xend174_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(105) & zeropad3D_D_CP_7327_elements(108) & zeropad3D_D_CP_7327_elements(111);
      gj_zeropad3D_D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	102 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	116 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2717/merge_stmt_2916_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_2717/merge_stmt_2916_PhiAck/$entry
      -- 
    zeropad3D_D_CP_7327_elements(113) <= OrReduce(zeropad3D_D_CP_7327_elements(102) & zeropad3D_D_CP_7327_elements(112));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	117 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2717/merge_stmt_2916_PhiAck/phi_stmt_2917_ack
      -- 
    phi_stmt_2917_ack_8687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2917_ack_0, ack => zeropad3D_D_CP_7327_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2717/merge_stmt_2916_PhiAck/phi_stmt_2923_ack
      -- 
    phi_stmt_2923_ack_8688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2923_ack_0, ack => zeropad3D_D_CP_7327_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	113 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2717/merge_stmt_2916_PhiAck/phi_stmt_2929_ack
      -- 
    phi_stmt_2929_ack_8689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2929_ack_0, ack => zeropad3D_D_CP_7327_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  place  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	114 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	23 
    -- CP-element group 117: 	24 
    -- CP-element group 117:  members (10) 
      -- CP-element group 117: 	 branch_block_stmt_2717/merge_stmt_2916_PhiAck/$exit
      -- CP-element group 117: 	 branch_block_stmt_2717/merge_stmt_2916__exit__
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948__entry__
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/$entry
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_update_start_
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_2717/assign_stmt_2941_to_assign_stmt_2948/type_cast_2940_Update/cr
      -- 
    rr_7750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(117), ack => type_cast_2940_inst_req_0); -- 
    cr_7755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(117), ack => type_cast_2940_inst_req_1); -- 
    zeropad3D_D_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(114) & zeropad3D_D_CP_7327_elements(115) & zeropad3D_D_CP_7327_elements(116);
      gj_zeropad3D_D_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  merge  fork  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	25 
    -- CP-element group 118: 	31 
    -- CP-element group 118: 	34 
    -- CP-element group 118: 	40 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	49 
    -- CP-element group 118: 	51 
    -- CP-element group 118: 	53 
    -- CP-element group 118: 	41 
    -- CP-element group 118: 	42 
    -- CP-element group 118: 	43 
    -- CP-element group 118: 	44 
    -- CP-element group 118: 	47 
    -- CP-element group 118:  members (33) 
      -- CP-element group 118: 	 branch_block_stmt_2717/merge_stmt_3032_PhiReqMerge
      -- CP-element group 118: 	 branch_block_stmt_2717/merge_stmt_3032__exit__
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088__entry__
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_update_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3036_Update/cr
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_update_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3041_Update/cr
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_update_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/type_cast_3075_Update/cr
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_update_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_update_start
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/array_obj_ref_3081_final_index_sum_regn_Update/req
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_complete/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/addr_of_3082_complete/req
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_update_start_
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/word_access_complete/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/word_access_complete/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/assign_stmt_3037_to_assign_stmt_3088/ptr_deref_3085_Update/word_access_complete/word_0/cr
      -- CP-element group 118: 	 branch_block_stmt_2717/merge_stmt_3032_PhiAck/$entry
      -- CP-element group 118: 	 branch_block_stmt_2717/merge_stmt_3032_PhiAck/$exit
      -- CP-element group 118: 	 branch_block_stmt_2717/merge_stmt_3032_PhiAck/dummy
      -- 
    rr_7966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => type_cast_3036_inst_req_0); -- 
    cr_7971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => type_cast_3036_inst_req_1); -- 
    rr_7980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => type_cast_3041_inst_req_0); -- 
    cr_7985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => type_cast_3041_inst_req_1); -- 
    cr_7999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => type_cast_3075_inst_req_1); -- 
    req_8030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => array_obj_ref_3081_index_offset_req_1); -- 
    req_8045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => addr_of_3082_final_reg_req_1); -- 
    cr_8095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(118), ack => ptr_deref_3085_store_0_req_1); -- 
    zeropad3D_D_CP_7327_elements(118) <= OrReduce(zeropad3D_D_CP_7327_elements(25) & zeropad3D_D_CP_7327_elements(31) & zeropad3D_D_CP_7327_elements(34) & zeropad3D_D_CP_7327_elements(40));
    -- CP-element group 119:  merge  fork  transition  place  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	54 
    -- CP-element group 119: 	74 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: 	76 
    -- CP-element group 119:  members (13) 
      -- CP-element group 119: 	 branch_block_stmt_2717/merge_stmt_3197_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2717/merge_stmt_3197__exit__
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215__entry__
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_update_start_
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/type_cast_3201_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_2717/assign_stmt_3202_to_assign_stmt_3215/$entry
      -- CP-element group 119: 	 branch_block_stmt_2717/merge_stmt_3197_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_2717/merge_stmt_3197_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_2717/merge_stmt_3197_PhiAck/dummy
      -- 
    cr_8349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(119), ack => type_cast_3201_inst_req_1); -- 
    rr_8344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(119), ack => type_cast_3201_inst_req_0); -- 
    zeropad3D_D_CP_7327_elements(119) <= OrReduce(zeropad3D_D_CP_7327_elements(54) & zeropad3D_D_CP_7327_elements(74));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	92 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Sample/ra
      -- 
    ra_8809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3324_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	92 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/Update/ca
      -- 
    ca_8814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3324_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	127 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/$exit
      -- CP-element group 122: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/$exit
      -- CP-element group 122: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3324/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_req
      -- 
    phi_stmt_3319_req_8815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3319_req_8815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(122), ack => phi_stmt_3319_req_1); -- 
    zeropad3D_D_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(120) & zeropad3D_D_CP_7327_elements(121);
      gj_zeropad3D_D_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	92 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Sample/ra
      -- 
    ra_8832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3316_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	92 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/Update/ca
      -- 
    ca_8837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3316_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/$exit
      -- CP-element group 125: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/$exit
      -- CP-element group 125: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3316/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_req
      -- 
    phi_stmt_3313_req_8838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3313_req_8838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(125), ack => phi_stmt_3313_req_0); -- 
    zeropad3D_D_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(123) & zeropad3D_D_CP_7327_elements(124);
      gj_zeropad3D_D_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  output  delay-element  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	92 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3325/$exit
      -- CP-element group 126: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3329_konst_delay_trans
      -- CP-element group 126: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_req
      -- 
    phi_stmt_3325_req_8846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3325_req_8846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(126), ack => phi_stmt_3325_req_0); -- 
    -- Element group zeropad3D_D_CP_7327_elements(126) is a control-delay.
    cp_element_126_delay: control_delay_element  generic map(name => " 126_delay", delay_value => 1)  port map(req => zeropad3D_D_CP_7327_elements(92), ack => zeropad3D_D_CP_7327_elements(126), clk => clk, reset =>reset);
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	122 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	138 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2717/ifx_xelse144_ifx_xend174_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(122) & zeropad3D_D_CP_7327_elements(125) & zeropad3D_D_CP_7327_elements(126);
      gj_zeropad3D_D_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	77 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Sample/ra
      -- 
    ra_8866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3322_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	77 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/Update/ca
      -- 
    ca_8871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3322_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	137 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/$exit
      -- CP-element group 130: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/$exit
      -- CP-element group 130: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/$exit
      -- CP-element group 130: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_sources/type_cast_3322/SplitProtocol/$exit
      -- CP-element group 130: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3319/phi_stmt_3319_req
      -- 
    phi_stmt_3319_req_8872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3319_req_8872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(130), ack => phi_stmt_3319_req_0); -- 
    zeropad3D_D_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(128) & zeropad3D_D_CP_7327_elements(129);
      gj_zeropad3D_D_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	77 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Sample/ra
      -- 
    ra_8889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3318_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	77 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/Update/ca
      -- 
    ca_8894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3318_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(132)); -- 
    -- CP-element group 133:  join  transition  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	137 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/$exit
      -- CP-element group 133: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/$exit
      -- CP-element group 133: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/$exit
      -- CP-element group 133: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_sources/type_cast_3318/SplitProtocol/$exit
      -- CP-element group 133: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3313/phi_stmt_3313_req
      -- 
    phi_stmt_3313_req_8895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3313_req_8895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(133), ack => phi_stmt_3313_req_1); -- 
    zeropad3D_D_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(131) & zeropad3D_D_CP_7327_elements(132);
      gj_zeropad3D_D_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	77 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Sample/ra
      -- 
    ra_8912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3331_inst_ack_0, ack => zeropad3D_D_CP_7327_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	77 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/Update/ca
      -- 
    ca_8917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3331_inst_ack_1, ack => zeropad3D_D_CP_7327_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (5) 
      -- CP-element group 136: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/$exit
      -- CP-element group 136: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/$exit
      -- CP-element group 136: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/$exit
      -- CP-element group 136: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_sources/type_cast_3331/SplitProtocol/$exit
      -- CP-element group 136: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/phi_stmt_3325/phi_stmt_3325_req
      -- 
    phi_stmt_3325_req_8918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3325_req_8918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_7327_elements(136), ack => phi_stmt_3325_req_1); -- 
    zeropad3D_D_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(134) & zeropad3D_D_CP_7327_elements(135);
      gj_zeropad3D_D_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	130 
    -- CP-element group 137: 	133 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_2717/ifx_xthen139_ifx_xend174_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(130) & zeropad3D_D_CP_7327_elements(133) & zeropad3D_D_CP_7327_elements(136);
      gj_zeropad3D_D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  merge  fork  transition  place  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	127 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	140 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_2717/merge_stmt_3312_PhiReqMerge
      -- CP-element group 138: 	 branch_block_stmt_2717/merge_stmt_3312_PhiAck/$entry
      -- 
    zeropad3D_D_CP_7327_elements(138) <= OrReduce(zeropad3D_D_CP_7327_elements(127) & zeropad3D_D_CP_7327_elements(137));
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_2717/merge_stmt_3312_PhiAck/phi_stmt_3313_ack
      -- 
    phi_stmt_3313_ack_8923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3313_ack_0, ack => zeropad3D_D_CP_7327_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_2717/merge_stmt_3312_PhiAck/phi_stmt_3319_ack
      -- 
    phi_stmt_3319_ack_8924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3319_ack_0, ack => zeropad3D_D_CP_7327_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_2717/merge_stmt_3312_PhiAck/phi_stmt_3325_ack
      -- 
    phi_stmt_3325_ack_8925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3325_ack_0, ack => zeropad3D_D_CP_7327_elements(141)); -- 
    -- CP-element group 142:  join  transition  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: 	140 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	1 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_2717/merge_stmt_3312_PhiAck/$exit
      -- 
    zeropad3D_D_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_7327_elements(139) & zeropad3D_D_CP_7327_elements(140) & zeropad3D_D_CP_7327_elements(141);
      gj_zeropad3D_D_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_7327_elements(142), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2817_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2832_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2847_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2871_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2886_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2912_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3069_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3152_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3177_wire : std_logic_vector(31 downto 0);
    signal LOAD_pad_2767_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2767_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom124_3163_resized : std_logic_vector(13 downto 0);
    signal R_idxprom124_3163_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom129_3188_resized : std_logic_vector(13 downto 0);
    signal R_idxprom129_3188_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3080_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3080_scaled : std_logic_vector(13 downto 0);
    signal add105_3125 : std_logic_vector(31 downto 0);
    signal add115_3140 : std_logic_vector(31 downto 0);
    signal add121_3145 : std_logic_vector(31 downto 0);
    signal add134_3208 : std_logic_vector(31 downto 0);
    signal add142_3228 : std_logic_vector(15 downto 0);
    signal add151_3258 : std_logic_vector(31 downto 0);
    signal add165_3300 : std_logic_vector(31 downto 0);
    signal add67_3020 : std_logic_vector(31 downto 0);
    signal add78_3057 : std_logic_vector(31 downto 0);
    signal add84_3062 : std_logic_vector(31 downto 0);
    signal add96_3120 : std_logic_vector(31 downto 0);
    signal add_2972 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3081_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3081_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3081_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3081_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3081_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3081_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3164_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3164_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3164_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3164_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3164_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3164_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3189_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3189_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3189_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3189_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3189_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3189_root_address : std_logic_vector(13 downto 0);
    signal arrayidx125_3166 : std_logic_vector(31 downto 0);
    signal arrayidx130_3191 : std_logic_vector(31 downto 0);
    signal arrayidx_3083 : std_logic_vector(31 downto 0);
    signal call_2720 : std_logic_vector(15 downto 0);
    signal cmp137_3215 : std_logic_vector(0 downto 0);
    signal cmp152_3263 : std_logic_vector(0 downto 0);
    signal cmp166_3305 : std_logic_vector(0 downto 0);
    signal cmp52_2977 : std_logic_vector(0 downto 0);
    signal cmp59_2996 : std_logic_vector(0 downto 0);
    signal cmp68_3025 : std_logic_vector(0 downto 0);
    signal cmp_2948 : std_logic_vector(0 downto 0);
    signal conv133_3202 : std_logic_vector(31 downto 0);
    signal conv136_2888 : std_logic_vector(31 downto 0);
    signal conv147_3241 : std_logic_vector(31 downto 0);
    signal conv160_3283 : std_logic_vector(31 downto 0);
    signal conv30_2819 : std_logic_vector(31 downto 0);
    signal conv34_2834 : std_logic_vector(31 downto 0);
    signal conv36_2849 : std_logic_vector(31 downto 0);
    signal conv43_2941 : std_logic_vector(31 downto 0);
    signal conv45_2858 : std_logic_vector(31 downto 0);
    signal conv4_2765 : std_logic_vector(15 downto 0);
    signal conv56_2989 : std_logic_vector(31 downto 0);
    signal conv72_3037 : std_logic_vector(31 downto 0);
    signal conv76_3042 : std_logic_vector(31 downto 0);
    signal conv80_2873 : std_logic_vector(31 downto 0);
    signal conv88_3095 : std_logic_vector(31 downto 0);
    signal conv98_2914 : std_logic_vector(31 downto 0);
    signal conv_2743 : std_logic_vector(15 downto 0);
    signal div3_2761 : std_logic_vector(31 downto 0);
    signal div_2739 : std_logic_vector(31 downto 0);
    signal iNsTr_11_2963 : std_logic_vector(31 downto 0);
    signal iNsTr_16_3249 : std_logic_vector(31 downto 0);
    signal iNsTr_17_3291 : std_logic_vector(31 downto 0);
    signal iNsTr_19_3011 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2729 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2751 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2776 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2788 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2800 : std_logic_vector(31 downto 0);
    signal idxprom124_3159 : std_logic_vector(63 downto 0);
    signal idxprom129_3184 : std_logic_vector(63 downto 0);
    signal idxprom_3076 : std_logic_vector(63 downto 0);
    signal inc157_3267 : std_logic_vector(15 downto 0);
    signal inc157x_xix_x2_3272 : std_logic_vector(15 downto 0);
    signal inc_3236 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_3313 : std_logic_vector(15 downto 0);
    signal ix_x2_2917 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_3319 : std_logic_vector(15 downto 0);
    signal jx_x1_2923 : std_logic_vector(15 downto 0);
    signal jx_x2_3278 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_3325 : std_logic_vector(15 downto 0);
    signal kx_x1_2929 : std_logic_vector(15 downto 0);
    signal mul104_3115 : std_logic_vector(31 downto 0);
    signal mul114_3130 : std_logic_vector(31 downto 0);
    signal mul120_3135 : std_logic_vector(31 downto 0);
    signal mul37_2854 : std_logic_vector(31 downto 0);
    signal mul77_3047 : std_logic_vector(31 downto 0);
    signal mul83_3052 : std_logic_vector(31 downto 0);
    signal mul95_3105 : std_logic_vector(31 downto 0);
    signal mul_2900 : std_logic_vector(31 downto 0);
    signal ptr_deref_2732_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2732_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2732_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2732_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2732_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2754_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2754_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2754_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2754_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2754_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2779_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2779_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2779_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2779_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2779_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2791_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2803_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2803_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2803_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2803_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2803_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2966_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2966_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2966_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2966_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2966_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3014_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3014_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3014_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3014_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3014_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3085_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3085_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3085_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3085_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3085_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3085_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3169_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3169_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3169_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3169_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3169_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3193_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3193_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3193_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3193_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3193_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3193_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3252_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3252_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3252_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3252_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3252_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3294_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3294_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3294_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3294_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3294_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext176_2840 : std_logic_vector(31 downto 0);
    signal sext177_2905 : std_logic_vector(31 downto 0);
    signal sext183_2825 : std_logic_vector(31 downto 0);
    signal sext184_2864 : std_logic_vector(31 downto 0);
    signal sext185_2879 : std_logic_vector(31 downto 0);
    signal sext_2810 : std_logic_vector(31 downto 0);
    signal shl_2894 : std_logic_vector(31 downto 0);
    signal shr123_3154 : std_logic_vector(31 downto 0);
    signal shr128_3179 : std_logic_vector(31 downto 0);
    signal shr_3071 : std_logic_vector(31 downto 0);
    signal sub103_3110 : std_logic_vector(31 downto 0);
    signal sub_3100 : std_logic_vector(31 downto 0);
    signal tmp126_3170 : std_logic_vector(63 downto 0);
    signal tmp148_3253 : std_logic_vector(31 downto 0);
    signal tmp161_3295 : std_logic_vector(31 downto 0);
    signal tmp18_2792 : std_logic_vector(31 downto 0);
    signal tmp21_2804 : std_logic_vector(31 downto 0);
    signal tmp2_2755 : std_logic_vector(31 downto 0);
    signal tmp49_2967 : std_logic_vector(31 downto 0);
    signal tmp64_3015 : std_logic_vector(31 downto 0);
    signal tmp6_2768 : std_logic_vector(7 downto 0);
    signal tmp9_2780 : std_logic_vector(31 downto 0);
    signal tmp_2733 : std_logic_vector(31 downto 0);
    signal type_cast_2737_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2759_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2808_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2813_wire : std_logic_vector(31 downto 0);
    signal type_cast_2816_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2823_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2828_wire : std_logic_vector(31 downto 0);
    signal type_cast_2831_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2843_wire : std_logic_vector(31 downto 0);
    signal type_cast_2846_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2862_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2867_wire : std_logic_vector(31 downto 0);
    signal type_cast_2870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2877_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2882_wire : std_logic_vector(31 downto 0);
    signal type_cast_2885_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2908_wire : std_logic_vector(31 downto 0);
    signal type_cast_2911_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2920_wire : std_logic_vector(15 downto 0);
    signal type_cast_2922_wire : std_logic_vector(15 downto 0);
    signal type_cast_2926_wire : std_logic_vector(15 downto 0);
    signal type_cast_2928_wire : std_logic_vector(15 downto 0);
    signal type_cast_2933_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2935_wire : std_logic_vector(15 downto 0);
    signal type_cast_2939_wire : std_logic_vector(31 downto 0);
    signal type_cast_2944_wire : std_logic_vector(31 downto 0);
    signal type_cast_2946_wire : std_logic_vector(31 downto 0);
    signal type_cast_2987_wire : std_logic_vector(31 downto 0);
    signal type_cast_2992_wire : std_logic_vector(31 downto 0);
    signal type_cast_2994_wire : std_logic_vector(31 downto 0);
    signal type_cast_3035_wire : std_logic_vector(31 downto 0);
    signal type_cast_3040_wire : std_logic_vector(31 downto 0);
    signal type_cast_3065_wire : std_logic_vector(31 downto 0);
    signal type_cast_3068_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3074_wire : std_logic_vector(63 downto 0);
    signal type_cast_3087_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3093_wire : std_logic_vector(31 downto 0);
    signal type_cast_3148_wire : std_logic_vector(31 downto 0);
    signal type_cast_3151_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3157_wire : std_logic_vector(63 downto 0);
    signal type_cast_3173_wire : std_logic_vector(31 downto 0);
    signal type_cast_3176_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3182_wire : std_logic_vector(63 downto 0);
    signal type_cast_3200_wire : std_logic_vector(31 downto 0);
    signal type_cast_3206_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3211_wire : std_logic_vector(31 downto 0);
    signal type_cast_3213_wire : std_logic_vector(31 downto 0);
    signal type_cast_3226_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3234_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3239_wire : std_logic_vector(31 downto 0);
    signal type_cast_3281_wire : std_logic_vector(31 downto 0);
    signal type_cast_3316_wire : std_logic_vector(15 downto 0);
    signal type_cast_3318_wire : std_logic_vector(15 downto 0);
    signal type_cast_3322_wire : std_logic_vector(15 downto 0);
    signal type_cast_3324_wire : std_logic_vector(15 downto 0);
    signal type_cast_3329_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3331_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_pad_2767_word_address_0 <= "0";
    array_obj_ref_3081_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3081_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3081_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3081_resized_base_address <= "00000000000000";
    array_obj_ref_3164_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3164_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3164_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3164_resized_base_address <= "00000000000000";
    array_obj_ref_3189_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3189_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3189_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3189_resized_base_address <= "00000000000000";
    iNsTr_11_2963 <= "00000000000000000000000000000011";
    iNsTr_16_3249 <= "00000000000000000000000000000100";
    iNsTr_17_3291 <= "00000000000000000000000000000011";
    iNsTr_19_3011 <= "00000000000000000000000000000100";
    iNsTr_2_2729 <= "00000000000000000000000000000100";
    iNsTr_3_2751 <= "00000000000000000000000000000011";
    iNsTr_4_2776 <= "00000000000000000000000000000101";
    iNsTr_5_2788 <= "00000000000000000000000000000101";
    iNsTr_6_2800 <= "00000000000000000000000000000100";
    ptr_deref_2732_word_offset_0 <= "0000000";
    ptr_deref_2754_word_offset_0 <= "0000000";
    ptr_deref_2779_word_offset_0 <= "0000000";
    ptr_deref_2791_word_offset_0 <= "0000000";
    ptr_deref_2803_word_offset_0 <= "0000000";
    ptr_deref_2966_word_offset_0 <= "0000000";
    ptr_deref_3014_word_offset_0 <= "0000000";
    ptr_deref_3085_word_offset_0 <= "00000000000000";
    ptr_deref_3169_word_offset_0 <= "00000000000000";
    ptr_deref_3193_word_offset_0 <= "00000000000000";
    ptr_deref_3252_word_offset_0 <= "0000000";
    ptr_deref_3294_word_offset_0 <= "0000000";
    type_cast_2737_wire_constant <= "00000000000000000000000000000001";
    type_cast_2759_wire_constant <= "00000000000000000000000000000001";
    type_cast_2808_wire_constant <= "00000000000000000000000000010000";
    type_cast_2816_wire_constant <= "00000000000000000000000000010000";
    type_cast_2823_wire_constant <= "00000000000000000000000000010000";
    type_cast_2831_wire_constant <= "00000000000000000000000000010000";
    type_cast_2838_wire_constant <= "00000000000000000000000000010000";
    type_cast_2846_wire_constant <= "00000000000000000000000000010000";
    type_cast_2862_wire_constant <= "00000000000000000000000000010000";
    type_cast_2870_wire_constant <= "00000000000000000000000000010000";
    type_cast_2877_wire_constant <= "00000000000000000000000000010000";
    type_cast_2885_wire_constant <= "00000000000000000000000000010000";
    type_cast_2892_wire_constant <= "00000000000000000000000000000001";
    type_cast_2898_wire_constant <= "00000000000000000000000000010000";
    type_cast_2911_wire_constant <= "00000000000000000000000000010000";
    type_cast_2933_wire_constant <= "0000000000000000";
    type_cast_3068_wire_constant <= "00000000000000000000000000000010";
    type_cast_3087_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3151_wire_constant <= "00000000000000000000000000000010";
    type_cast_3176_wire_constant <= "00000000000000000000000000000010";
    type_cast_3206_wire_constant <= "00000000000000000000000000000100";
    type_cast_3226_wire_constant <= "0000000000000100";
    type_cast_3234_wire_constant <= "0000000000000001";
    type_cast_3329_wire_constant <= "0000000000000000";
    phi_stmt_2917: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2920_wire & type_cast_2922_wire;
      req <= phi_stmt_2917_req_0 & phi_stmt_2917_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2917",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2917_ack_0,
          idata => idata,
          odata => ix_x2_2917,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2917
    phi_stmt_2923: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2926_wire & type_cast_2928_wire;
      req <= phi_stmt_2923_req_0 & phi_stmt_2923_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2923",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2923_ack_0,
          idata => idata,
          odata => jx_x1_2923,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2923
    phi_stmt_2929: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2933_wire_constant & type_cast_2935_wire;
      req <= phi_stmt_2929_req_0 & phi_stmt_2929_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2929",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2929_ack_0,
          idata => idata,
          odata => kx_x1_2929,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2929
    phi_stmt_3313: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3316_wire & type_cast_3318_wire;
      req <= phi_stmt_3313_req_0 & phi_stmt_3313_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3313",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3313_ack_0,
          idata => idata,
          odata => ix_x1x_xph_3313,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3313
    phi_stmt_3319: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3322_wire & type_cast_3324_wire;
      req <= phi_stmt_3319_req_0 & phi_stmt_3319_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3319",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3319_ack_0,
          idata => idata,
          odata => jx_x0x_xph_3319,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3319
    phi_stmt_3325: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3329_wire_constant & type_cast_3331_wire;
      req <= phi_stmt_3325_req_0 & phi_stmt_3325_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3325",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3325_ack_0,
          idata => idata,
          odata => kx_x0x_xph_3325,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3325
    -- flow-through select operator MUX_3277_inst
    jx_x2_3278 <= conv_2743 when (cmp152_3263(0) /=  '0') else inc_3236;
    addr_of_3082_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3082_final_reg_req_0;
      addr_of_3082_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3082_final_reg_req_1;
      addr_of_3082_final_reg_ack_1<= rack(0);
      addr_of_3082_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3082_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3081_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3083,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3165_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3165_final_reg_req_0;
      addr_of_3165_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3165_final_reg_req_1;
      addr_of_3165_final_reg_ack_1<= rack(0);
      addr_of_3165_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3165_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3164_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx125_3166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3190_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3190_final_reg_req_0;
      addr_of_3190_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3190_final_reg_req_1;
      addr_of_3190_final_reg_ack_1<= rack(0);
      addr_of_3190_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3190_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3189_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx130_3191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2742_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2742_inst_req_0;
      type_cast_2742_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2742_inst_req_1;
      type_cast_2742_inst_ack_1<= rack(0);
      type_cast_2742_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2742_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2739,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2764_inst_req_0;
      type_cast_2764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2764_inst_req_1;
      type_cast_2764_inst_ack_1<= rack(0);
      type_cast_2764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div3_2761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2813_inst
    process(sext_2810) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2810(31 downto 0);
      type_cast_2813_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2818_inst
    process(ASHR_i32_i32_2817_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2817_wire(31 downto 0);
      conv30_2819 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2828_inst
    process(sext183_2825) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext183_2825(31 downto 0);
      type_cast_2828_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2833_inst
    process(ASHR_i32_i32_2832_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2832_wire(31 downto 0);
      conv34_2834 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2843_inst
    process(sext176_2840) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext176_2840(31 downto 0);
      type_cast_2843_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2848_inst
    process(ASHR_i32_i32_2847_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2847_wire(31 downto 0);
      conv36_2849 <= tmp_var; -- 
    end process;
    type_cast_2857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2857_inst_req_0;
      type_cast_2857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2857_inst_req_1;
      type_cast_2857_inst_ack_1<= rack(0);
      type_cast_2857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6_2768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_2858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2867_inst
    process(sext184_2864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext184_2864(31 downto 0);
      type_cast_2867_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2872_inst
    process(ASHR_i32_i32_2871_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2871_wire(31 downto 0);
      conv80_2873 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2882_inst
    process(sext185_2879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext185_2879(31 downto 0);
      type_cast_2882_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2887_inst
    process(ASHR_i32_i32_2886_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2886_wire(31 downto 0);
      conv136_2888 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2908_inst
    process(sext177_2905) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext177_2905(31 downto 0);
      type_cast_2908_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2913_inst
    process(ASHR_i32_i32_2912_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2912_wire(31 downto 0);
      conv98_2914 <= tmp_var; -- 
    end process;
    type_cast_2920_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2920_inst_req_0;
      type_cast_2920_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2920_inst_req_1;
      type_cast_2920_inst_ack_1<= rack(0);
      type_cast_2920_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2920_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_2765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2920_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2922_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2922_inst_req_0;
      type_cast_2922_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2922_inst_req_1;
      type_cast_2922_inst_ack_1<= rack(0);
      type_cast_2922_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2922_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_3313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2922_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2926_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2926_inst_req_0;
      type_cast_2926_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2926_inst_req_1;
      type_cast_2926_inst_ack_1<= rack(0);
      type_cast_2926_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2926_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2926_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2928_inst_req_0;
      type_cast_2928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2928_inst_req_1;
      type_cast_2928_inst_ack_1<= rack(0);
      type_cast_2928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_3319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2928_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2935_inst_req_0;
      type_cast_2935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2935_inst_req_1;
      type_cast_2935_inst_ack_1<= rack(0);
      type_cast_2935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_3325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2935_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2940_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2940_inst_req_0;
      type_cast_2940_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2940_inst_req_1;
      type_cast_2940_inst_ack_1<= rack(0);
      type_cast_2940_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2940_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2939_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_2941,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2944_inst
    process(conv43_2941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv43_2941(31 downto 0);
      type_cast_2944_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2946_inst
    process(conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv45_2858(31 downto 0);
      type_cast_2946_wire <= tmp_var; -- 
    end process;
    type_cast_2988_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2988_inst_req_0;
      type_cast_2988_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2988_inst_req_1;
      type_cast_2988_inst_ack_1<= rack(0);
      type_cast_2988_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2988_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2987_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_2989,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2992_inst
    process(conv56_2989) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv56_2989(31 downto 0);
      type_cast_2992_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2994_inst
    process(conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv45_2858(31 downto 0);
      type_cast_2994_wire <= tmp_var; -- 
    end process;
    type_cast_3036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3036_inst_req_0;
      type_cast_3036_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3036_inst_req_1;
      type_cast_3036_inst_ack_1<= rack(0);
      type_cast_3036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3036_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3035_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_3037,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3041_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3041_inst_req_0;
      type_cast_3041_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3041_inst_req_1;
      type_cast_3041_inst_ack_1<= rack(0);
      type_cast_3041_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3041_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3040_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_3042,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3065_inst
    process(add84_3062) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add84_3062(31 downto 0);
      type_cast_3065_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3070_inst
    process(ASHR_i32_i32_3069_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3069_wire(31 downto 0);
      shr_3071 <= tmp_var; -- 
    end process;
    type_cast_3075_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3075_inst_req_0;
      type_cast_3075_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3075_inst_req_1;
      type_cast_3075_inst_ack_1<= rack(0);
      type_cast_3075_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3075_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3074_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3076,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3094_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3094_inst_req_0;
      type_cast_3094_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3094_inst_req_1;
      type_cast_3094_inst_ack_1<= rack(0);
      type_cast_3094_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3094_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3093_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3148_inst
    process(add105_3125) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add105_3125(31 downto 0);
      type_cast_3148_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3153_inst
    process(ASHR_i32_i32_3152_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3152_wire(31 downto 0);
      shr123_3154 <= tmp_var; -- 
    end process;
    type_cast_3158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3158_inst_req_0;
      type_cast_3158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3158_inst_req_1;
      type_cast_3158_inst_ack_1<= rack(0);
      type_cast_3158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3157_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom124_3159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3173_inst
    process(add121_3145) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add121_3145(31 downto 0);
      type_cast_3173_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3178_inst
    process(ASHR_i32_i32_3177_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3177_wire(31 downto 0);
      shr128_3179 <= tmp_var; -- 
    end process;
    type_cast_3183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3183_inst_req_0;
      type_cast_3183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3183_inst_req_1;
      type_cast_3183_inst_ack_1<= rack(0);
      type_cast_3183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3182_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom129_3184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3201_inst_req_0;
      type_cast_3201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3201_inst_req_1;
      type_cast_3201_inst_ack_1<= rack(0);
      type_cast_3201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3200_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv133_3202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3211_inst
    process(add134_3208) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add134_3208(31 downto 0);
      type_cast_3211_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3213_inst
    process(conv136_2888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv136_2888(31 downto 0);
      type_cast_3213_wire <= tmp_var; -- 
    end process;
    type_cast_3240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3240_inst_req_0;
      type_cast_3240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3240_inst_req_1;
      type_cast_3240_inst_ack_1<= rack(0);
      type_cast_3240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3239_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_3241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3266_inst_req_0;
      type_cast_3266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3266_inst_req_1;
      type_cast_3266_inst_ack_1<= rack(0);
      type_cast_3266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp152_3263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc157_3267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3282_inst_req_0;
      type_cast_3282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3282_inst_req_1;
      type_cast_3282_inst_ack_1<= rack(0);
      type_cast_3282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3281_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_3283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3316_inst_req_0;
      type_cast_3316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3316_inst_req_1;
      type_cast_3316_inst_ack_1<= rack(0);
      type_cast_3316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc157x_xix_x2_3272,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3316_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3318_inst_req_0;
      type_cast_3318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3318_inst_req_1;
      type_cast_3318_inst_ack_1<= rack(0);
      type_cast_3318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_2917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3318_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3322_inst_req_0;
      type_cast_3322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3322_inst_req_1;
      type_cast_3322_inst_ack_1<= rack(0);
      type_cast_3322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_2923,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3322_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3324_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3324_inst_req_0;
      type_cast_3324_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3324_inst_req_1;
      type_cast_3324_inst_ack_1<= rack(0);
      type_cast_3324_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3324_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_3278,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3324_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3331_inst_req_0;
      type_cast_3331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3331_inst_req_1;
      type_cast_3331_inst_ack_1<= rack(0);
      type_cast_3331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add142_3228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3331_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_pad_2767_gather_scatter
    process(LOAD_pad_2767_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2767_data_0;
      ov(7 downto 0) := iv;
      tmp6_2768 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3081_index_1_rename
    process(R_idxprom_3080_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3080_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3080_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3081_index_1_resize
    process(idxprom_3076) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3076;
      ov := iv(13 downto 0);
      R_idxprom_3080_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3081_root_address_inst
    process(array_obj_ref_3081_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3081_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3081_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3164_index_1_rename
    process(R_idxprom124_3163_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom124_3163_resized;
      ov(13 downto 0) := iv;
      R_idxprom124_3163_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3164_index_1_resize
    process(idxprom124_3159) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom124_3159;
      ov := iv(13 downto 0);
      R_idxprom124_3163_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3164_root_address_inst
    process(array_obj_ref_3164_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3164_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3164_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3189_index_1_rename
    process(R_idxprom129_3188_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom129_3188_resized;
      ov(13 downto 0) := iv;
      R_idxprom129_3188_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3189_index_1_resize
    process(idxprom129_3184) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom129_3184;
      ov := iv(13 downto 0);
      R_idxprom129_3188_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3189_root_address_inst
    process(array_obj_ref_3189_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3189_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3189_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2732_addr_0
    process(ptr_deref_2732_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2732_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2732_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2732_base_resize
    process(iNsTr_2_2729) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2729;
      ov := iv(6 downto 0);
      ptr_deref_2732_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2732_gather_scatter
    process(ptr_deref_2732_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2732_data_0;
      ov(31 downto 0) := iv;
      tmp_2733 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2732_root_address_inst
    process(ptr_deref_2732_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2732_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2732_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_addr_0
    process(ptr_deref_2754_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2754_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2754_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_base_resize
    process(iNsTr_3_2751) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2751;
      ov := iv(6 downto 0);
      ptr_deref_2754_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_gather_scatter
    process(ptr_deref_2754_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2754_data_0;
      ov(31 downto 0) := iv;
      tmp2_2755 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_root_address_inst
    process(ptr_deref_2754_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2754_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2754_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2779_addr_0
    process(ptr_deref_2779_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2779_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2779_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2779_base_resize
    process(iNsTr_4_2776) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2776;
      ov := iv(6 downto 0);
      ptr_deref_2779_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2779_gather_scatter
    process(ptr_deref_2779_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2779_data_0;
      ov(31 downto 0) := iv;
      tmp9_2780 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2779_root_address_inst
    process(ptr_deref_2779_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2779_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2779_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_addr_0
    process(ptr_deref_2791_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2791_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2791_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_base_resize
    process(iNsTr_5_2788) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2788;
      ov := iv(6 downto 0);
      ptr_deref_2791_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_gather_scatter
    process(ptr_deref_2791_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2791_data_0;
      ov(31 downto 0) := iv;
      tmp18_2792 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_root_address_inst
    process(ptr_deref_2791_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2791_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2791_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2803_addr_0
    process(ptr_deref_2803_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2803_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2803_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2803_base_resize
    process(iNsTr_6_2800) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2800;
      ov := iv(6 downto 0);
      ptr_deref_2803_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2803_gather_scatter
    process(ptr_deref_2803_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2803_data_0;
      ov(31 downto 0) := iv;
      tmp21_2804 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2803_root_address_inst
    process(ptr_deref_2803_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2803_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2803_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2966_addr_0
    process(ptr_deref_2966_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2966_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2966_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2966_base_resize
    process(iNsTr_11_2963) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_11_2963;
      ov := iv(6 downto 0);
      ptr_deref_2966_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2966_gather_scatter
    process(ptr_deref_2966_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2966_data_0;
      ov(31 downto 0) := iv;
      tmp49_2967 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2966_root_address_inst
    process(ptr_deref_2966_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2966_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2966_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3014_addr_0
    process(ptr_deref_3014_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3014_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3014_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3014_base_resize
    process(iNsTr_19_3011) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_19_3011;
      ov := iv(6 downto 0);
      ptr_deref_3014_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3014_gather_scatter
    process(ptr_deref_3014_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3014_data_0;
      ov(31 downto 0) := iv;
      tmp64_3015 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3014_root_address_inst
    process(ptr_deref_3014_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3014_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3014_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3085_addr_0
    process(ptr_deref_3085_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3085_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3085_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3085_base_resize
    process(arrayidx_3083) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3083;
      ov := iv(13 downto 0);
      ptr_deref_3085_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3085_gather_scatter
    process(type_cast_3087_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3087_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3085_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3085_root_address_inst
    process(ptr_deref_3085_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3085_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3085_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3169_addr_0
    process(ptr_deref_3169_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3169_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3169_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3169_base_resize
    process(arrayidx125_3166) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx125_3166;
      ov := iv(13 downto 0);
      ptr_deref_3169_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3169_gather_scatter
    process(ptr_deref_3169_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3169_data_0;
      ov(63 downto 0) := iv;
      tmp126_3170 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3169_root_address_inst
    process(ptr_deref_3169_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3169_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3169_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3193_addr_0
    process(ptr_deref_3193_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3193_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3193_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3193_base_resize
    process(arrayidx130_3191) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx130_3191;
      ov := iv(13 downto 0);
      ptr_deref_3193_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3193_gather_scatter
    process(tmp126_3170) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp126_3170;
      ov(63 downto 0) := iv;
      ptr_deref_3193_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3193_root_address_inst
    process(ptr_deref_3193_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3193_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3193_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3252_addr_0
    process(ptr_deref_3252_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3252_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3252_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3252_base_resize
    process(iNsTr_16_3249) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_16_3249;
      ov := iv(6 downto 0);
      ptr_deref_3252_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3252_gather_scatter
    process(ptr_deref_3252_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3252_data_0;
      ov(31 downto 0) := iv;
      tmp148_3253 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3252_root_address_inst
    process(ptr_deref_3252_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3252_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3252_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3294_addr_0
    process(ptr_deref_3294_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3294_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3294_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3294_base_resize
    process(iNsTr_17_3291) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_3291;
      ov := iv(6 downto 0);
      ptr_deref_3294_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3294_gather_scatter
    process(ptr_deref_3294_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3294_data_0;
      ov(31 downto 0) := iv;
      tmp161_3295 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3294_root_address_inst
    process(ptr_deref_3294_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3294_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3294_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_2949_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2948;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2949_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2949_branch_req_0,
          ack0 => if_stmt_2949_branch_ack_0,
          ack1 => if_stmt_2949_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2978_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp52_2977;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2978_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2978_branch_req_0,
          ack0 => if_stmt_2978_branch_ack_0,
          ack1 => if_stmt_2978_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2997_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp59_2996;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2997_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2997_branch_req_0,
          ack0 => if_stmt_2997_branch_ack_0,
          ack1 => if_stmt_2997_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3026_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_3025;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3026_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3026_branch_req_0,
          ack0 => if_stmt_3026_branch_ack_0,
          ack1 => if_stmt_3026_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3216_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp137_3215;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3216_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3216_branch_req_0,
          ack0 => if_stmt_3216_branch_ack_0,
          ack1 => if_stmt_3216_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3306_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp166_3305;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3306_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3306_branch_req_0,
          ack0 => if_stmt_3306_branch_ack_0,
          ack1 => if_stmt_3306_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3227_inst
    process(kx_x1_2929) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_2929, type_cast_3226_wire_constant, tmp_var);
      add142_3228 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3235_inst
    process(jx_x1_2923) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_2923, type_cast_3234_wire_constant, tmp_var);
      inc_3236 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3271_inst
    process(inc157_3267, ix_x2_2917) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc157_3267, ix_x2_2917, tmp_var);
      inc157x_xix_x2_3272 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2971_inst
    process(tmp49_2967, conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp49_2967, conv45_2858, tmp_var);
      add_2972 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3019_inst
    process(tmp64_3015, conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp64_3015, conv45_2858, tmp_var);
      add67_3020 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3056_inst
    process(mul77_3047, mul83_3052) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul77_3047, mul83_3052, tmp_var);
      add78_3057 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3061_inst
    process(add78_3057, conv72_3037) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add78_3057, conv72_3037, tmp_var);
      add84_3062 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3119_inst
    process(conv88_3095, mul104_3115) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv88_3095, mul104_3115, tmp_var);
      add96_3120 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3124_inst
    process(add96_3120, mul95_3105) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add96_3120, mul95_3105, tmp_var);
      add105_3125 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3139_inst
    process(mul114_3130, mul120_3135) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul114_3130, mul120_3135, tmp_var);
      add115_3140 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3144_inst
    process(add115_3140, conv88_3095) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add115_3140, conv88_3095, tmp_var);
      add121_3145 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3207_inst
    process(conv133_3202) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv133_3202, type_cast_3206_wire_constant, tmp_var);
      add134_3208 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3257_inst
    process(tmp148_3253, shl_2894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp148_3253, shl_2894, tmp_var);
      add151_3258 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3299_inst
    process(tmp161_3295, shl_2894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp161_3295, shl_2894, tmp_var);
      add165_3300 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2817_inst
    process(type_cast_2813_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2813_wire, type_cast_2816_wire_constant, tmp_var);
      ASHR_i32_i32_2817_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2832_inst
    process(type_cast_2828_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2828_wire, type_cast_2831_wire_constant, tmp_var);
      ASHR_i32_i32_2832_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2847_inst
    process(type_cast_2843_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2843_wire, type_cast_2846_wire_constant, tmp_var);
      ASHR_i32_i32_2847_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2871_inst
    process(type_cast_2867_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2867_wire, type_cast_2870_wire_constant, tmp_var);
      ASHR_i32_i32_2871_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2886_inst
    process(type_cast_2882_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2882_wire, type_cast_2885_wire_constant, tmp_var);
      ASHR_i32_i32_2886_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2912_inst
    process(type_cast_2908_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2908_wire, type_cast_2911_wire_constant, tmp_var);
      ASHR_i32_i32_2912_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3069_inst
    process(type_cast_3065_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3065_wire, type_cast_3068_wire_constant, tmp_var);
      ASHR_i32_i32_3069_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3152_inst
    process(type_cast_3148_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3148_wire, type_cast_3151_wire_constant, tmp_var);
      ASHR_i32_i32_3152_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3177_inst
    process(type_cast_3173_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3173_wire, type_cast_3176_wire_constant, tmp_var);
      ASHR_i32_i32_3177_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3262_inst
    process(conv147_3241, add151_3258) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv147_3241, add151_3258, tmp_var);
      cmp152_3263 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3304_inst
    process(conv160_3283, add165_3300) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv160_3283, add165_3300, tmp_var);
      cmp166_3305 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2738_inst
    process(tmp_2733) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2733, type_cast_2737_wire_constant, tmp_var);
      div_2739 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2760_inst
    process(tmp2_2755) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2755, type_cast_2759_wire_constant, tmp_var);
      div3_2761 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2853_inst
    process(conv36_2849, conv34_2834) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv36_2849, conv34_2834, tmp_var);
      mul37_2854 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2904_inst
    process(mul_2900, conv30_2819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_2900, conv30_2819, tmp_var);
      sext177_2905 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3046_inst
    process(conv76_3042, conv34_2834) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv76_3042, conv34_2834, tmp_var);
      mul77_3047 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3051_inst
    process(conv43_2941, conv80_2873) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv43_2941, conv80_2873, tmp_var);
      mul83_3052 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3104_inst
    process(sub_3100, conv136_2888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_3100, conv136_2888, tmp_var);
      mul95_3105 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3114_inst
    process(sub103_3110, conv98_2914) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub103_3110, conv98_2914, tmp_var);
      mul104_3115 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3129_inst
    process(conv56_2989, conv34_2834) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv56_2989, conv34_2834, tmp_var);
      mul114_3130 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3134_inst
    process(conv43_2941, conv80_2873) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv43_2941, conv80_2873, tmp_var);
      mul120_3135 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2809_inst
    process(tmp_2733) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp_2733, type_cast_2808_wire_constant, tmp_var);
      sext_2810 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2824_inst
    process(tmp18_2792) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp18_2792, type_cast_2823_wire_constant, tmp_var);
      sext183_2825 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2839_inst
    process(tmp21_2804) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp21_2804, type_cast_2838_wire_constant, tmp_var);
      sext176_2840 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2863_inst
    process(mul37_2854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul37_2854, type_cast_2862_wire_constant, tmp_var);
      sext184_2864 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2878_inst
    process(tmp9_2780) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp9_2780, type_cast_2877_wire_constant, tmp_var);
      sext185_2879 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2893_inst
    process(conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv45_2858, type_cast_2892_wire_constant, tmp_var);
      shl_2894 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2899_inst
    process(tmp9_2780) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp9_2780, type_cast_2898_wire_constant, tmp_var);
      mul_2900 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2947_inst
    process(type_cast_2944_wire, type_cast_2946_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2944_wire, type_cast_2946_wire, tmp_var);
      cmp_2948 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2995_inst
    process(type_cast_2992_wire, type_cast_2994_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2992_wire, type_cast_2994_wire, tmp_var);
      cmp59_2996 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3214_inst
    process(type_cast_3211_wire, type_cast_3213_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3211_wire, type_cast_3213_wire, tmp_var);
      cmp137_3215 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3099_inst
    process(conv56_2989, conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv56_2989, conv45_2858, tmp_var);
      sub_3100 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3109_inst
    process(conv43_2941, conv45_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv43_2941, conv45_2858, tmp_var);
      sub103_3110 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2976_inst
    process(conv43_2941, add_2972) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv43_2941, add_2972, tmp_var);
      cmp52_2977 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3024_inst
    process(conv56_2989, add67_3020) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv56_2989, add67_3020, tmp_var);
      cmp68_3025 <= tmp_var; --
    end process;
    -- shared split operator group (49) : array_obj_ref_3081_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3080_scaled;
      array_obj_ref_3081_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3081_index_offset_req_0;
      array_obj_ref_3081_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3081_index_offset_req_1;
      array_obj_ref_3081_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : array_obj_ref_3164_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom124_3163_scaled;
      array_obj_ref_3164_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3164_index_offset_req_0;
      array_obj_ref_3164_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3164_index_offset_req_1;
      array_obj_ref_3164_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : array_obj_ref_3189_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom129_3188_scaled;
      array_obj_ref_3189_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3189_index_offset_req_0;
      array_obj_ref_3189_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3189_index_offset_req_1;
      array_obj_ref_3189_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- unary operator type_cast_2939_inst
    process(ix_x2_2917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_2917, tmp_var);
      type_cast_2939_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2987_inst
    process(jx_x1_2923) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2923, tmp_var);
      type_cast_2987_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3035_inst
    process(kx_x1_2929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2929, tmp_var);
      type_cast_3035_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3040_inst
    process(jx_x1_2923) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2923, tmp_var);
      type_cast_3040_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3074_inst
    process(shr_3071) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3071, tmp_var);
      type_cast_3074_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3093_inst
    process(kx_x1_2929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2929, tmp_var);
      type_cast_3093_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3157_inst
    process(shr123_3154) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr123_3154, tmp_var);
      type_cast_3157_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3182_inst
    process(shr128_3179) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr128_3179, tmp_var);
      type_cast_3182_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3200_inst
    process(kx_x1_2929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2929, tmp_var);
      type_cast_3200_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3239_inst
    process(inc_3236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3236, tmp_var);
      type_cast_3239_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3281_inst
    process(inc157x_xix_x2_3272) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc157x_xix_x2_3272, tmp_var);
      type_cast_3281_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_pad_2767_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_pad_2767_load_0_req_0;
      LOAD_pad_2767_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_pad_2767_load_0_req_1;
      LOAD_pad_2767_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_2767_word_address_0;
      LOAD_pad_2767_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(0 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2966_load_0 ptr_deref_2779_load_0 ptr_deref_2754_load_0 ptr_deref_2732_load_0 ptr_deref_3294_load_0 ptr_deref_3252_load_0 ptr_deref_3014_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(48 downto 0);
      signal data_out: std_logic_vector(223 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= ptr_deref_2966_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_2779_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_2754_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2732_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3294_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_3252_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3014_load_0_req_0;
      ptr_deref_2966_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_2779_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_2754_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2732_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3294_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_3252_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3014_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= ptr_deref_2966_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_2779_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_2754_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2732_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3294_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_3252_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3014_load_0_req_1;
      ptr_deref_2966_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_2779_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_2754_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2732_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3294_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_3252_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3014_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2966_word_address_0 & ptr_deref_2779_word_address_0 & ptr_deref_2754_word_address_0 & ptr_deref_2732_word_address_0 & ptr_deref_3294_word_address_0 & ptr_deref_3252_word_address_0 & ptr_deref_3014_word_address_0;
      ptr_deref_2966_data_0 <= data_out(223 downto 192);
      ptr_deref_2779_data_0 <= data_out(191 downto 160);
      ptr_deref_2754_data_0 <= data_out(159 downto 128);
      ptr_deref_2732_data_0 <= data_out(127 downto 96);
      ptr_deref_3294_data_0 <= data_out(95 downto 64);
      ptr_deref_3252_data_0 <= data_out(63 downto 32);
      ptr_deref_3014_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 7,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 7,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2791_load_0 ptr_deref_2803_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2791_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2803_load_0_req_0;
      ptr_deref_2791_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2803_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2791_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2803_load_0_req_1;
      ptr_deref_2791_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2803_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2791_word_address_0 & ptr_deref_2803_word_address_0;
      ptr_deref_2791_data_0 <= data_out(63 downto 32);
      ptr_deref_2803_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(6 downto 0),
          mtag => memory_space_4_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_3169_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3169_load_0_req_0;
      ptr_deref_3169_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3169_load_0_req_1;
      ptr_deref_3169_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3169_word_address_0;
      ptr_deref_3169_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_3085_store_0 ptr_deref_3193_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3085_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3193_store_0_req_0;
      ptr_deref_3085_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3193_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3085_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3193_store_0_req_1;
      ptr_deref_3085_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3193_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3085_word_address_0 & ptr_deref_3193_word_address_0;
      data_in <= ptr_deref_3085_data_0 & ptr_deref_3193_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_starting_2719_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_starting_2719_inst_req_0;
      RPIPE_Block3_starting_2719_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_starting_2719_inst_req_1;
      RPIPE_Block3_starting_2719_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2720 <= data_out(15 downto 0);
      Block3_starting_read_0_gI: SplitGuardInterface generic map(name => "Block3_starting_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block3_starting_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_starting_pipe_read_req(0),
          oack => Block3_starting_pipe_read_ack(0),
          odata => Block3_starting_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_complete_3336_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_complete_3336_inst_req_0;
      WPIPE_Block3_complete_3336_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_complete_3336_inst_req_1;
      WPIPE_Block3_complete_3336_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2720;
      Block3_complete_write_0_gI: SplitGuardInterface generic map(name => "Block3_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_complete", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_complete_pipe_write_req(0),
          oack => Block3_complete_pipe_write_ack(0),
          odata => Block3_complete_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(79 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(7 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(99 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_complete_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      Block2_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_starting_pipe_write_data : out  std_logic_vector(15 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- declarations related to module zeropad3D_A
  component zeropad3D_A is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_A
  signal zeropad3D_A_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_A_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_A_start_req : std_logic;
  signal zeropad3D_A_start_ack : std_logic;
  signal zeropad3D_A_fin_req   : std_logic;
  signal zeropad3D_A_fin_ack : std_logic;
  -- declarations related to module zeropad3D_B
  component zeropad3D_B is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block1_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_B
  signal zeropad3D_B_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_B_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_B_start_req : std_logic;
  signal zeropad3D_B_start_ack : std_logic;
  signal zeropad3D_B_fin_req   : std_logic;
  signal zeropad3D_B_fin_ack : std_logic;
  -- declarations related to module zeropad3D_C
  component zeropad3D_C is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block2_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_C
  signal zeropad3D_C_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_C_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_C_start_req : std_logic;
  signal zeropad3D_C_start_ack : std_logic;
  signal zeropad3D_C_fin_req   : std_logic;
  signal zeropad3D_C_fin_ack : std_logic;
  -- declarations related to module zeropad3D_D
  component zeropad3D_D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block3_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_starting_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_complete_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_D
  signal zeropad3D_D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_D_start_req : std_logic;
  signal zeropad3D_D_start_ack : std_logic;
  signal zeropad3D_D_fin_req   : std_logic;
  signal zeropad3D_D_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_complete
  signal Block0_complete_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_complete
  signal Block0_complete_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_starting
  signal Block0_starting_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_starting
  signal Block0_starting_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_complete
  signal Block1_complete_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_complete
  signal Block1_complete_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_starting
  signal Block1_starting_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_starting
  signal Block1_starting_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_complete
  signal Block2_complete_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_complete
  signal Block2_complete_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_starting
  signal Block2_starting_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_starting
  signal Block2_starting_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_complete
  signal Block3_complete_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_complete
  signal Block3_complete_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_starting
  signal Block3_starting_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_starting
  signal Block3_starting_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(4 downto 4),
      memory_space_4_lr_ack => memory_space_4_lr_ack(4 downto 4),
      memory_space_4_lr_addr => memory_space_4_lr_addr(34 downto 28),
      memory_space_4_lr_tag => memory_space_4_lr_tag(99 downto 80),
      memory_space_4_lc_req => memory_space_4_lc_req(4 downto 4),
      memory_space_4_lc_ack => memory_space_4_lc_ack(4 downto 4),
      memory_space_4_lc_data => memory_space_4_lc_data(159 downto 128),
      memory_space_4_lc_tag => memory_space_4_lc_tag(9 downto 8),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(4 downto 4),
      memory_space_3_lr_ack => memory_space_3_lr_ack(4 downto 4),
      memory_space_3_lr_addr => memory_space_3_lr_addr(34 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(104 downto 84),
      memory_space_3_lc_req => memory_space_3_lc_req(4 downto 4),
      memory_space_3_lc_ack => memory_space_3_lc_ack(4 downto 4),
      memory_space_3_lc_data => memory_space_3_lc_data(159 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(14 downto 12),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(20 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(6 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(31 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(19 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(1 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(0 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(7 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(0 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      Block0_complete_pipe_read_req => Block0_complete_pipe_read_req(0 downto 0),
      Block0_complete_pipe_read_ack => Block0_complete_pipe_read_ack(0 downto 0),
      Block0_complete_pipe_read_data => Block0_complete_pipe_read_data(15 downto 0),
      Block1_complete_pipe_read_req => Block1_complete_pipe_read_req(0 downto 0),
      Block1_complete_pipe_read_ack => Block1_complete_pipe_read_ack(0 downto 0),
      Block1_complete_pipe_read_data => Block1_complete_pipe_read_data(15 downto 0),
      Block3_complete_pipe_read_req => Block3_complete_pipe_read_req(0 downto 0),
      Block3_complete_pipe_read_ack => Block3_complete_pipe_read_ack(0 downto 0),
      Block3_complete_pipe_read_data => Block3_complete_pipe_read_data(15 downto 0),
      Block2_complete_pipe_read_req => Block2_complete_pipe_read_req(0 downto 0),
      Block2_complete_pipe_read_ack => Block2_complete_pipe_read_ack(0 downto 0),
      Block2_complete_pipe_read_data => Block2_complete_pipe_read_data(15 downto 0),
      Block1_starting_pipe_write_req => Block1_starting_pipe_write_req(0 downto 0),
      Block1_starting_pipe_write_ack => Block1_starting_pipe_write_ack(0 downto 0),
      Block1_starting_pipe_write_data => Block1_starting_pipe_write_data(15 downto 0),
      Block0_starting_pipe_write_req => Block0_starting_pipe_write_req(0 downto 0),
      Block0_starting_pipe_write_ack => Block0_starting_pipe_write_ack(0 downto 0),
      Block0_starting_pipe_write_data => Block0_starting_pipe_write_data(15 downto 0),
      Block3_starting_pipe_write_req => Block3_starting_pipe_write_req(0 downto 0),
      Block3_starting_pipe_write_ack => Block3_starting_pipe_write_ack(0 downto 0),
      Block3_starting_pipe_write_data => Block3_starting_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      Block2_starting_pipe_write_req => Block2_starting_pipe_write_req(0 downto 0),
      Block2_starting_pipe_write_ack => Block2_starting_pipe_write_ack(0 downto 0),
      Block2_starting_pipe_write_data => Block2_starting_pipe_write_data(15 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  -- module zeropad3D_A
  zeropad3D_A_instance:zeropad3D_A-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_A_start_req,
      start_ack => zeropad3D_A_start_ack,
      fin_req => zeropad3D_A_fin_req,
      fin_ack => zeropad3D_A_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 21),
      memory_space_3_lr_tag => memory_space_3_lr_tag(83 downto 63),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 96),
      memory_space_3_lc_tag => memory_space_3_lc_tag(11 downto 9),
      memory_space_4_lr_req => memory_space_4_lr_req(3 downto 3),
      memory_space_4_lr_ack => memory_space_4_lr_ack(3 downto 3),
      memory_space_4_lr_addr => memory_space_4_lr_addr(27 downto 21),
      memory_space_4_lr_tag => memory_space_4_lr_tag(79 downto 60),
      memory_space_4_lc_req => memory_space_4_lc_req(3 downto 3),
      memory_space_4_lc_ack => memory_space_4_lc_ack(3 downto 3),
      memory_space_4_lc_data => memory_space_4_lc_data(127 downto 96),
      memory_space_4_lc_tag => memory_space_4_lc_tag(7 downto 6),
      memory_space_5_lr_req => memory_space_5_lr_req(3 downto 3),
      memory_space_5_lr_ack => memory_space_5_lr_ack(3 downto 3),
      memory_space_5_lr_addr => memory_space_5_lr_addr(3 downto 3),
      memory_space_5_lr_tag => memory_space_5_lr_tag(75 downto 57),
      memory_space_5_lc_req => memory_space_5_lc_req(3 downto 3),
      memory_space_5_lc_ack => memory_space_5_lc_ack(3 downto 3),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 24),
      memory_space_5_lc_tag => memory_space_5_lc_tag(3 downto 3),
      memory_space_0_sr_req => memory_space_0_sr_req(3 downto 3),
      memory_space_0_sr_ack => memory_space_0_sr_ack(3 downto 3),
      memory_space_0_sr_addr => memory_space_0_sr_addr(55 downto 42),
      memory_space_0_sr_data => memory_space_0_sr_data(255 downto 192),
      memory_space_0_sr_tag => memory_space_0_sr_tag(79 downto 60),
      memory_space_0_sc_req => memory_space_0_sc_req(3 downto 3),
      memory_space_0_sc_ack => memory_space_0_sc_ack(3 downto 3),
      memory_space_0_sc_tag => memory_space_0_sc_tag(7 downto 6),
      Block0_starting_pipe_read_req => Block0_starting_pipe_read_req(0 downto 0),
      Block0_starting_pipe_read_ack => Block0_starting_pipe_read_ack(0 downto 0),
      Block0_starting_pipe_read_data => Block0_starting_pipe_read_data(15 downto 0),
      Block0_complete_pipe_write_req => Block0_complete_pipe_write_req(0 downto 0),
      Block0_complete_pipe_write_ack => Block0_complete_pipe_write_ack(0 downto 0),
      Block0_complete_pipe_write_data => Block0_complete_pipe_write_data(15 downto 0),
      tag_in => zeropad3D_A_tag_in,
      tag_out => zeropad3D_A_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_A_tag_in <= (others => '0');
  zeropad3D_A_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_A_start_req, start_ack => zeropad3D_A_start_ack,  fin_req => zeropad3D_A_fin_req,  fin_ack => zeropad3D_A_fin_ack);
  -- module zeropad3D_B
  zeropad3D_B_instance:zeropad3D_B-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_B_start_req,
      start_ack => zeropad3D_B_start_ack,
      fin_req => zeropad3D_B_fin_req,
      fin_ack => zeropad3D_B_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(20 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(62 downto 42),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(95 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(8 downto 6),
      memory_space_4_lr_req => memory_space_4_lr_req(2 downto 2),
      memory_space_4_lr_ack => memory_space_4_lr_ack(2 downto 2),
      memory_space_4_lr_addr => memory_space_4_lr_addr(20 downto 14),
      memory_space_4_lr_tag => memory_space_4_lr_tag(59 downto 40),
      memory_space_4_lc_req => memory_space_4_lc_req(2 downto 2),
      memory_space_4_lc_ack => memory_space_4_lc_ack(2 downto 2),
      memory_space_4_lc_data => memory_space_4_lc_data(95 downto 64),
      memory_space_4_lc_tag => memory_space_4_lc_tag(5 downto 4),
      memory_space_5_lr_req => memory_space_5_lr_req(2 downto 2),
      memory_space_5_lr_ack => memory_space_5_lr_ack(2 downto 2),
      memory_space_5_lr_addr => memory_space_5_lr_addr(2 downto 2),
      memory_space_5_lr_tag => memory_space_5_lr_tag(56 downto 38),
      memory_space_5_lc_req => memory_space_5_lc_req(2 downto 2),
      memory_space_5_lc_ack => memory_space_5_lc_ack(2 downto 2),
      memory_space_5_lc_data => memory_space_5_lc_data(23 downto 16),
      memory_space_5_lc_tag => memory_space_5_lc_tag(2 downto 2),
      memory_space_0_sr_req => memory_space_0_sr_req(2 downto 2),
      memory_space_0_sr_ack => memory_space_0_sr_ack(2 downto 2),
      memory_space_0_sr_addr => memory_space_0_sr_addr(41 downto 28),
      memory_space_0_sr_data => memory_space_0_sr_data(191 downto 128),
      memory_space_0_sr_tag => memory_space_0_sr_tag(59 downto 40),
      memory_space_0_sc_req => memory_space_0_sc_req(2 downto 2),
      memory_space_0_sc_ack => memory_space_0_sc_ack(2 downto 2),
      memory_space_0_sc_tag => memory_space_0_sc_tag(5 downto 4),
      Block1_starting_pipe_read_req => Block1_starting_pipe_read_req(0 downto 0),
      Block1_starting_pipe_read_ack => Block1_starting_pipe_read_ack(0 downto 0),
      Block1_starting_pipe_read_data => Block1_starting_pipe_read_data(15 downto 0),
      Block1_complete_pipe_write_req => Block1_complete_pipe_write_req(0 downto 0),
      Block1_complete_pipe_write_ack => Block1_complete_pipe_write_ack(0 downto 0),
      Block1_complete_pipe_write_data => Block1_complete_pipe_write_data(15 downto 0),
      tag_in => zeropad3D_B_tag_in,
      tag_out => zeropad3D_B_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_B_tag_in <= (others => '0');
  zeropad3D_B_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_B_start_req, start_ack => zeropad3D_B_start_ack,  fin_req => zeropad3D_B_fin_req,  fin_ack => zeropad3D_B_fin_ack);
  -- module zeropad3D_C
  zeropad3D_C_instance:zeropad3D_C-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_C_start_req,
      start_ack => zeropad3D_C_start_ack,
      fin_req => zeropad3D_C_fin_req,
      fin_ack => zeropad3D_C_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(41 downto 21),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(5 downto 3),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(13 downto 7),
      memory_space_4_lr_tag => memory_space_4_lr_tag(39 downto 20),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(63 downto 32),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 2),
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(1 downto 1),
      memory_space_5_lr_tag => memory_space_5_lr_tag(37 downto 19),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(15 downto 8),
      memory_space_5_lc_tag => memory_space_5_lc_tag(1 downto 1),
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(27 downto 14),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      Block2_starting_pipe_read_req => Block2_starting_pipe_read_req(0 downto 0),
      Block2_starting_pipe_read_ack => Block2_starting_pipe_read_ack(0 downto 0),
      Block2_starting_pipe_read_data => Block2_starting_pipe_read_data(15 downto 0),
      Block2_complete_pipe_write_req => Block2_complete_pipe_write_req(0 downto 0),
      Block2_complete_pipe_write_ack => Block2_complete_pipe_write_ack(0 downto 0),
      Block2_complete_pipe_write_data => Block2_complete_pipe_write_data(15 downto 0),
      tag_in => zeropad3D_C_tag_in,
      tag_out => zeropad3D_C_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_C_tag_in <= (others => '0');
  zeropad3D_C_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_C_start_req, start_ack => zeropad3D_C_start_ack,  fin_req => zeropad3D_C_fin_req,  fin_ack => zeropad3D_C_fin_ack);
  -- module zeropad3D_D
  zeropad3D_D_instance:zeropad3D_D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_D_start_req,
      start_ack => zeropad3D_D_start_ack,
      fin_req => zeropad3D_D_fin_req,
      fin_ack => zeropad3D_D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(20 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(6 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(19 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(1 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(0 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(7 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Block3_starting_pipe_read_req => Block3_starting_pipe_read_req(0 downto 0),
      Block3_starting_pipe_read_ack => Block3_starting_pipe_read_ack(0 downto 0),
      Block3_starting_pipe_read_data => Block3_starting_pipe_read_data(15 downto 0),
      Block3_complete_pipe_write_req => Block3_complete_pipe_write_req(0 downto 0),
      Block3_complete_pipe_write_ack => Block3_complete_pipe_write_ack(0 downto 0),
      Block3_complete_pipe_write_data => Block3_complete_pipe_write_data(15 downto 0),
      tag_in => zeropad3D_D_tag_in,
      tag_out => zeropad3D_D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_D_tag_in <= (others => '0');
  zeropad3D_D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_D_start_req, start_ack => zeropad3D_D_start_ack,  fin_req => zeropad3D_D_fin_req,  fin_ack => zeropad3D_D_fin_ack);
  Block0_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_complete_pipe_read_req,
      read_ack => Block0_complete_pipe_read_ack,
      read_data => Block0_complete_pipe_read_data,
      write_req => Block0_complete_pipe_write_req,
      write_ack => Block0_complete_pipe_write_ack,
      write_data => Block0_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_starting_pipe_read_req,
      read_ack => Block0_starting_pipe_read_ack,
      read_data => Block0_starting_pipe_read_data,
      write_req => Block0_starting_pipe_write_req,
      write_ack => Block0_starting_pipe_write_ack,
      write_data => Block0_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_complete_pipe_read_req,
      read_ack => Block1_complete_pipe_read_ack,
      read_data => Block1_complete_pipe_read_data,
      write_req => Block1_complete_pipe_write_req,
      write_ack => Block1_complete_pipe_write_ack,
      write_data => Block1_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_starting_pipe_read_req,
      read_ack => Block1_starting_pipe_read_ack,
      read_data => Block1_starting_pipe_read_data,
      write_req => Block1_starting_pipe_write_req,
      write_ack => Block1_starting_pipe_write_ack,
      write_data => Block1_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_complete_pipe_read_req,
      read_ack => Block2_complete_pipe_read_ack,
      read_data => Block2_complete_pipe_read_data,
      write_req => Block2_complete_pipe_write_req,
      write_ack => Block2_complete_pipe_write_ack,
      write_data => Block2_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_starting_pipe_read_req,
      read_ack => Block2_starting_pipe_read_ack,
      read_data => Block2_starting_pipe_read_data,
      write_req => Block2_starting_pipe_write_req,
      write_ack => Block2_starting_pipe_write_ack,
      write_data => Block2_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_complete_pipe_read_req,
      read_ack => Block3_complete_pipe_read_ack,
      read_data => Block3_complete_pipe_read_data,
      write_req => Block3_complete_pipe_write_req,
      write_ack => Block3_complete_pipe_write_ack,
      write_data => Block3_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_starting_pipe_read_req,
      read_ack => Block3_starting_pipe_read_ack,
      read_data => Block3_starting_pipe_read_data,
      write_req => Block3_starting_pipe_write_req,
      write_ack => Block3_starting_pipe_write_ack,
      write_data => Block3_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 4,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyROM_memory_space_2: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
