-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_3_start: Boolean;
  signal timer_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_15_load_0_req_0 : boolean;
  signal LOAD_count_15_load_0_ack_0 : boolean;
  signal LOAD_count_15_load_0_req_1 : boolean;
  signal LOAD_count_15_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_3: Block -- control-path 
    signal timer_CP_3_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_3_elements(0) <= timer_CP_3_start;
    timer_CP_3_symbol <= timer_CP_3_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_16/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_sample_start_
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_update_start_
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Update/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_16/LOAD_count_15_Update/word_access_complete/word_0/cr
      -- 
    cr_35_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_35_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_3_elements(0), ack => LOAD_count_15_load_0_req_1); -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_3_elements(0), ack => LOAD_count_15_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_16/LOAD_count_15_sample_completed_
      -- CP-element group 1: 	 assign_stmt_16/LOAD_count_15_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_16/LOAD_count_15_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_16/LOAD_count_15_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_16/LOAD_count_15_Sample/word_access_start/word_0/ra
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_15_load_0_ack_0, ack => timer_CP_3_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_16/$exit
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/LOAD_count_15_Merge/merge_ack
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_update_completed_
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/$exit
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/LOAD_count_15_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/LOAD_count_15_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_16/LOAD_count_15_Update/LOAD_count_15_Merge/merge_req
      -- 
    ca_36_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_15_load_0_ack_1, ack => timer_CP_3_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_15_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_15_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_15_word_address_0 <= "0";
    -- equivalence LOAD_count_15_gather_scatter
    process(LOAD_count_15_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_15_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_15_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_15_load_0_req_0;
      LOAD_count_15_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_15_load_0_req_1;
      LOAD_count_15_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_15_word_address_0;
      LOAD_count_15_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_42_start: Boolean;
  signal timerDaemon_CP_42_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_20_branch_req_0 : boolean;
  signal phi_stmt_22_req_1 : boolean;
  signal phi_stmt_22_req_0 : boolean;
  signal phi_stmt_22_ack_0 : boolean;
  signal ADD_u64_u64_28_inst_req_0 : boolean;
  signal ADD_u64_u64_28_inst_ack_0 : boolean;
  signal ADD_u64_u64_28_inst_req_1 : boolean;
  signal ADD_u64_u64_28_inst_ack_1 : boolean;
  signal STORE_count_30_store_0_req_0 : boolean;
  signal STORE_count_30_store_0_ack_0 : boolean;
  signal STORE_count_30_store_0_req_1 : boolean;
  signal STORE_count_30_store_0_ack_1 : boolean;
  signal do_while_stmt_20_branch_ack_0 : boolean;
  signal do_while_stmt_20_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_42_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_42_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_42_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_42_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_42: Block -- control-path 
    signal timerDaemon_CP_42_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_42_elements(0) <= timerDaemon_CP_42_start;
    timerDaemon_CP_42_symbol <= timerDaemon_CP_42_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_19/$entry
      -- CP-element group 0: 	 branch_block_stmt_19/branch_block_stmt_19__entry__
      -- CP-element group 0: 	 branch_block_stmt_19/do_while_stmt_20__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_19/$exit
      -- CP-element group 1: 	 branch_block_stmt_19/branch_block_stmt_19__exit__
      -- CP-element group 1: 	 branch_block_stmt_19/do_while_stmt_20__exit__
      -- 
    timerDaemon_CP_42_elements(1) <= timerDaemon_CP_42_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_19/do_while_stmt_20/$entry
      -- CP-element group 2: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20__entry__
      -- 
    timerDaemon_CP_42_elements(2) <= timerDaemon_CP_42_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20__exit__
      -- 
    -- Element group timerDaemon_CP_42_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_19/do_while_stmt_20/loop_back
      -- 
    -- Element group timerDaemon_CP_42_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_19/do_while_stmt_20/condition_done
      -- CP-element group 5: 	 branch_block_stmt_19/do_while_stmt_20/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_19/do_while_stmt_20/loop_taken/$entry
      -- 
    timerDaemon_CP_42_elements(5) <= timerDaemon_CP_42_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_19/do_while_stmt_20/loop_body_done
      -- 
    timerDaemon_CP_42_elements(6) <= timerDaemon_CP_42_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_42_elements(7) <= timerDaemon_CP_42_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_42_elements(8) <= timerDaemon_CP_42_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_42_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/condition_evaluated
      -- 
    condition_evaluated_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(10), ack => do_while_stmt_20_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(15) & timerDaemon_CP_42_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(12) & timerDaemon_CP_42_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(9) & timerDaemon_CP_42_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_start_
      -- CP-element group 13: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(9) & timerDaemon_CP_42_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_42_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_42_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_loopback_trigger
      -- 
    timerDaemon_CP_42_elements(16) <= timerDaemon_CP_42_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_loopback_sample_req_ps
      -- 
    phi_stmt_22_loopback_sample_req_81_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_22_loopback_sample_req_81_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(17), ack => phi_stmt_22_req_1); -- 
    -- Element group timerDaemon_CP_42_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_entry_trigger
      -- 
    timerDaemon_CP_42_elements(18) <= timerDaemon_CP_42_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_entry_sample_req_ps
      -- 
    phi_stmt_22_entry_sample_req_84_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_22_entry_sample_req_84_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(19), ack => phi_stmt_22_req_0); -- 
    -- Element group timerDaemon_CP_42_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_phi_mux_ack_ps
      -- 
    phi_stmt_22_phi_mux_ack_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_22_ack_0, ack => timerDaemon_CP_42_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_completed_
      -- 
    -- Element group timerDaemon_CP_42_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_start_
      -- 
    -- Element group timerDaemon_CP_42_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_completed__ps
      -- 
    timerDaemon_CP_42_elements(23) <= timerDaemon_CP_42_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_completed_
      -- 
    -- Element group timerDaemon_CP_42_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_42_elements(22), ack => timerDaemon_CP_42_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_42_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_update_start__ps
      -- 
    -- Element group timerDaemon_CP_42_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Sample/rr
      -- 
    rr_108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(27), ack => ADD_u64_u64_28_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(25) & timerDaemon_CP_42_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_update_start_
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Update/cr
      -- 
    cr_113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(28), ack => ADD_u64_u64_28_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(26) & timerDaemon_CP_42_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Sample/ra
      -- 
    ra_109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_28_inst_ack_0, ack => timerDaemon_CP_42_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u64_u64_28_Update/ca
      -- 
    ca_114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_28_inst_ack_1, ack => timerDaemon_CP_42_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/STORE_count_30_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/STORE_count_30_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/STORE_count_30_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/STORE_count_30_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/word_access_start/word_0/rr
      -- 
    rr_136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(31), ack => STORE_count_30_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(9) & timerDaemon_CP_42_elements(15) & timerDaemon_CP_42_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_update_start_
      -- CP-element group 32: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/word_access_complete/word_0/cr
      -- 
    cr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_42_elements(32), ack => STORE_count_30_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_42_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Sample/word_access_start/word_0/ra
      -- 
    ra_137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_30_store_0_ack_0, ack => timerDaemon_CP_42_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/STORE_count_30_Update/word_access_complete/word_0/ca
      -- 
    ca_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_30_store_0_ack_1, ack => timerDaemon_CP_42_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_42_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_42_elements(9), ack => timerDaemon_CP_42_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_42_elements(14) & timerDaemon_CP_42_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_42_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_19/do_while_stmt_20/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_19/do_while_stmt_20/loop_exit/ack
      -- 
    ack_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_20_branch_ack_0, ack => timerDaemon_CP_42_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_19/do_while_stmt_20/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_19/do_while_stmt_20/loop_taken/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_20_branch_ack_1, ack => timerDaemon_CP_42_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_19/do_while_stmt_20/$exit
      -- 
    timerDaemon_CP_42_elements(39) <= timerDaemon_CP_42_elements(3);
    timerDaemon_do_while_stmt_20_terminator_158: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_20_terminator_158", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_42_elements(6),loop_continue => timerDaemon_CP_42_elements(38),loop_terminate => timerDaemon_CP_42_elements(37),loop_back => timerDaemon_CP_42_elements(4),loop_exit => timerDaemon_CP_42_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_22_phi_seq_115_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_42_elements(18);
      timerDaemon_CP_42_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_42_elements(21);
      timerDaemon_CP_42_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_42_elements(23);
      timerDaemon_CP_42_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_42_elements(16);
      timerDaemon_CP_42_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_42_elements(29);
      timerDaemon_CP_42_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_42_elements(30);
      timerDaemon_CP_42_elements(17) <= phi_mux_reqs(1);
      phi_stmt_22_phi_seq_115 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_22_phi_seq_115") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_42_elements(11), 
          phi_sample_ack => timerDaemon_CP_42_elements(14), 
          phi_update_req => timerDaemon_CP_42_elements(13), 
          phi_update_ack => timerDaemon_CP_42_elements(15), 
          phi_mux_ack => timerDaemon_CP_42_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_67_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_42_elements(7);
        preds(1)  <= timerDaemon_CP_42_elements(8);
        entry_tmerge_67 : transition_merge -- 
          generic map(name => " entry_tmerge_67")
          port map (preds => preds, symbol_out => timerDaemon_CP_42_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_28_wire : std_logic_vector(63 downto 0);
    signal STORE_count_30_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_30_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_27_wire_constant : std_logic_vector(63 downto 0);
    signal konst_34_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_22 : std_logic_vector(63 downto 0);
    signal type_cast_25_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_30_word_address_0 <= "0";
    konst_27_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_34_wire_constant <= "1";
    type_cast_25_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_22: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_25_wire_constant & ADD_u64_u64_28_wire;
      req <= phi_stmt_22_req_0 & phi_stmt_22_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_22",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_22_ack_0,
          idata => idata,
          odata => ncount_22,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_22
    -- equivalence STORE_count_30_gather_scatter
    process(ncount_22) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_22;
      ov(63 downto 0) := iv;
      STORE_count_30_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_20_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_34_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_20_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_20_branch_req_0,
          ack0 => do_while_stmt_20_branch_ack_0,
          ack1 => do_while_stmt_20_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_28_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_22;
      ADD_u64_u64_28_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_28_inst_req_0;
      ADD_u64_u64_28_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_28_inst_req_1;
      ADD_u64_u64_28_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_30_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_30_store_0_req_0;
      STORE_count_30_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_30_store_0_req_1;
      STORE_count_30_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_30_word_address_0;
      data_in <= STORE_count_30_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad_same is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad_same;
architecture zeropad_same_arch of zeropad_same is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad_same_CP_159_start: Boolean;
  signal zeropad_same_CP_159_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal next_input_dim2_740_588_buf_ack_0 : boolean;
  signal phi_stmt_585_ack_0 : boolean;
  signal array_obj_ref_956_index_offset_req_0 : boolean;
  signal next_input_dim2_740_588_buf_req_1 : boolean;
  signal next_input_dim2_740_588_buf_ack_1 : boolean;
  signal type_cast_787_inst_ack_0 : boolean;
  signal addr_of_515_final_reg_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_881_inst_req_0 : boolean;
  signal next_input_dim0_756_580_buf_ack_0 : boolean;
  signal next_input_dim0_756_580_buf_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_890_inst_ack_0 : boolean;
  signal addr_of_515_final_reg_ack_0 : boolean;
  signal phi_stmt_577_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_881_inst_ack_0 : boolean;
  signal phi_stmt_581_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_878_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_878_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_878_inst_req_0 : boolean;
  signal type_cast_837_inst_req_0 : boolean;
  signal next_input_dim1_750_584_buf_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_887_inst_req_1 : boolean;
  signal next_input_dim1_750_584_buf_req_1 : boolean;
  signal type_cast_787_inst_ack_1 : boolean;
  signal type_cast_58_inst_req_0 : boolean;
  signal type_cast_58_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_890_inst_req_1 : boolean;
  signal type_cast_58_inst_req_1 : boolean;
  signal type_cast_58_inst_ack_1 : boolean;
  signal addr_of_515_final_reg_req_0 : boolean;
  signal type_cast_807_inst_ack_1 : boolean;
  signal phi_stmt_585_req_1 : boolean;
  signal if_stmt_458_branch_req_0 : boolean;
  signal next_input_dim2_740_588_buf_req_0 : boolean;
  signal type_cast_787_inst_req_1 : boolean;
  signal addr_of_957_final_reg_ack_0 : boolean;
  signal phi_stmt_585_req_0 : boolean;
  signal if_stmt_458_branch_ack_0 : boolean;
  signal if_stmt_458_branch_ack_1 : boolean;
  signal addr_of_515_final_reg_ack_1 : boolean;
  signal type_cast_797_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_878_inst_ack_1 : boolean;
  signal type_cast_45_inst_req_0 : boolean;
  signal type_cast_45_inst_ack_0 : boolean;
  signal type_cast_45_inst_req_1 : boolean;
  signal type_cast_45_inst_ack_1 : boolean;
  signal phi_stmt_577_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_ack_0 : boolean;
  signal addr_of_957_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_ack_1 : boolean;
  signal next_input_dim1_750_584_buf_ack_0 : boolean;
  signal next_input_dim1_750_584_buf_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_884_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_884_inst_ack_1 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 : boolean;
  signal if_stmt_533_branch_req_0 : boolean;
  signal array_obj_ref_514_index_offset_ack_0 : boolean;
  signal type_cast_70_inst_req_0 : boolean;
  signal type_cast_70_inst_ack_0 : boolean;
  signal type_cast_70_inst_req_1 : boolean;
  signal type_cast_70_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_ack_1 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal call_stmt_777_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_881_inst_ack_1 : boolean;
  signal array_obj_ref_514_index_offset_ack_1 : boolean;
  signal phi_stmt_581_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_0 : boolean;
  signal type_cast_837_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 : boolean;
  signal array_obj_ref_514_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal addr_of_957_final_reg_ack_1 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal call_stmt_544_call_ack_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal phi_stmt_577_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_req_1 : boolean;
  signal call_stmt_544_call_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_ack_1 : boolean;
  signal type_cast_782_inst_ack_0 : boolean;
  signal type_cast_837_inst_ack_0 : boolean;
  signal type_cast_797_inst_req_1 : boolean;
  signal type_cast_108_inst_req_0 : boolean;
  signal type_cast_108_inst_ack_0 : boolean;
  signal type_cast_108_inst_req_1 : boolean;
  signal type_cast_108_inst_ack_1 : boolean;
  signal array_obj_ref_514_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_1 : boolean;
  signal call_stmt_544_call_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 : boolean;
  signal next_input_dim0_756_580_buf_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_887_inst_ack_1 : boolean;
  signal type_cast_120_inst_req_0 : boolean;
  signal call_stmt_544_call_req_0 : boolean;
  signal type_cast_120_inst_ack_0 : boolean;
  signal type_cast_120_inst_req_1 : boolean;
  signal type_cast_120_inst_ack_1 : boolean;
  signal array_obj_ref_956_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_ack_1 : boolean;
  signal ptr_deref_518_store_0_ack_1 : boolean;
  signal type_cast_133_inst_req_0 : boolean;
  signal type_cast_133_inst_ack_0 : boolean;
  signal type_cast_133_inst_req_1 : boolean;
  signal type_cast_133_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 : boolean;
  signal call_stmt_777_call_req_1 : boolean;
  signal next_input_dim0_756_580_buf_req_1 : boolean;
  signal ptr_deref_518_store_0_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_884_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_890_inst_ack_1 : boolean;
  signal type_cast_145_inst_req_0 : boolean;
  signal type_cast_145_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_1 : boolean;
  signal type_cast_797_inst_ack_0 : boolean;
  signal type_cast_145_inst_ack_1 : boolean;
  signal type_cast_782_inst_ack_1 : boolean;
  signal do_while_stmt_575_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_ack_0 : boolean;
  signal phi_stmt_581_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_ack_1 : boolean;
  signal type_cast_158_inst_req_0 : boolean;
  signal type_cast_158_inst_ack_0 : boolean;
  signal type_cast_158_inst_req_1 : boolean;
  signal type_cast_158_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_881_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 : boolean;
  signal type_cast_782_inst_req_1 : boolean;
  signal type_cast_170_inst_req_0 : boolean;
  signal type_cast_170_inst_ack_0 : boolean;
  signal type_cast_170_inst_req_1 : boolean;
  signal type_cast_170_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_884_inst_ack_0 : boolean;
  signal type_cast_183_inst_req_0 : boolean;
  signal type_cast_183_inst_ack_0 : boolean;
  signal type_cast_183_inst_req_1 : boolean;
  signal type_cast_183_inst_ack_1 : boolean;
  signal ptr_deref_518_store_0_ack_0 : boolean;
  signal type_cast_193_inst_req_0 : boolean;
  signal type_cast_193_inst_ack_0 : boolean;
  signal type_cast_193_inst_req_1 : boolean;
  signal if_stmt_533_branch_ack_0 : boolean;
  signal type_cast_193_inst_ack_1 : boolean;
  signal ptr_deref_518_store_0_req_0 : boolean;
  signal type_cast_202_inst_req_0 : boolean;
  signal type_cast_202_inst_ack_0 : boolean;
  signal type_cast_202_inst_req_1 : boolean;
  signal type_cast_202_inst_ack_1 : boolean;
  signal type_cast_485_inst_ack_1 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_485_inst_req_1 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_837_inst_ack_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal type_cast_782_inst_req_0 : boolean;
  signal type_cast_220_inst_req_0 : boolean;
  signal if_stmt_533_branch_ack_1 : boolean;
  signal type_cast_220_inst_ack_0 : boolean;
  signal type_cast_220_inst_req_1 : boolean;
  signal type_cast_220_inst_ack_1 : boolean;
  signal type_cast_485_inst_ack_0 : boolean;
  signal type_cast_485_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_890_inst_req_0 : boolean;
  signal if_stmt_234_branch_req_0 : boolean;
  signal if_stmt_234_branch_ack_1 : boolean;
  signal if_stmt_234_branch_ack_0 : boolean;
  signal type_cast_265_inst_req_0 : boolean;
  signal type_cast_265_inst_ack_0 : boolean;
  signal type_cast_265_inst_req_1 : boolean;
  signal type_cast_265_inst_ack_1 : boolean;
  signal array_obj_ref_294_index_offset_req_0 : boolean;
  signal array_obj_ref_294_index_offset_ack_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal array_obj_ref_294_index_offset_req_1 : boolean;
  signal array_obj_ref_294_index_offset_ack_1 : boolean;
  signal addr_of_295_final_reg_req_0 : boolean;
  signal addr_of_295_final_reg_ack_0 : boolean;
  signal addr_of_295_final_reg_req_1 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal addr_of_295_final_reg_ack_1 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal ptr_deref_961_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_1 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 : boolean;
  signal type_cast_302_inst_req_0 : boolean;
  signal type_cast_302_inst_ack_0 : boolean;
  signal type_cast_302_inst_req_1 : boolean;
  signal type_cast_302_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_ack_1 : boolean;
  signal type_cast_315_inst_req_0 : boolean;
  signal type_cast_315_inst_ack_0 : boolean;
  signal type_cast_315_inst_req_1 : boolean;
  signal type_cast_315_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 : boolean;
  signal type_cast_827_inst_req_0 : boolean;
  signal type_cast_827_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_887_inst_req_0 : boolean;
  signal type_cast_333_inst_req_0 : boolean;
  signal type_cast_333_inst_ack_0 : boolean;
  signal type_cast_333_inst_req_1 : boolean;
  signal type_cast_333_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal type_cast_827_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_887_inst_ack_0 : boolean;
  signal type_cast_351_inst_req_0 : boolean;
  signal type_cast_351_inst_ack_0 : boolean;
  signal type_cast_351_inst_req_1 : boolean;
  signal type_cast_351_inst_ack_1 : boolean;
  signal type_cast_797_inst_ack_1 : boolean;
  signal array_obj_ref_956_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_365_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_365_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_365_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_365_inst_ack_1 : boolean;
  signal type_cast_827_inst_ack_1 : boolean;
  signal if_stmt_900_branch_req_0 : boolean;
  signal type_cast_369_inst_req_0 : boolean;
  signal type_cast_369_inst_ack_0 : boolean;
  signal type_cast_369_inst_req_1 : boolean;
  signal type_cast_369_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_ack_1 : boolean;
  signal type_cast_387_inst_req_0 : boolean;
  signal type_cast_387_inst_ack_0 : boolean;
  signal type_cast_387_inst_req_1 : boolean;
  signal type_cast_387_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_401_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_401_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_401_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_401_inst_ack_1 : boolean;
  signal type_cast_405_inst_req_0 : boolean;
  signal type_cast_405_inst_ack_0 : boolean;
  signal type_cast_405_inst_req_1 : boolean;
  signal type_cast_405_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_ack_1 : boolean;
  signal type_cast_423_inst_req_0 : boolean;
  signal type_cast_423_inst_ack_0 : boolean;
  signal type_cast_423_inst_req_1 : boolean;
  signal type_cast_423_inst_ack_1 : boolean;
  signal ptr_deref_431_store_0_req_0 : boolean;
  signal ptr_deref_431_store_0_ack_0 : boolean;
  signal ptr_deref_431_store_0_req_1 : boolean;
  signal ptr_deref_431_store_0_ack_1 : boolean;
  signal if_stmt_445_branch_req_0 : boolean;
  signal if_stmt_445_branch_ack_1 : boolean;
  signal if_stmt_445_branch_ack_0 : boolean;
  signal type_cast_787_inst_req_0 : boolean;
  signal phi_stmt_589_req_1 : boolean;
  signal addr_of_957_final_reg_req_0 : boolean;
  signal phi_stmt_589_req_0 : boolean;
  signal phi_stmt_589_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_875_inst_ack_1 : boolean;
  signal add_dest_dim0_init_567_591_buf_req_0 : boolean;
  signal add_dest_dim0_init_567_591_buf_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_875_inst_req_1 : boolean;
  signal add_dest_dim0_init_567_591_buf_req_1 : boolean;
  signal add_dest_dim0_init_567_591_buf_ack_1 : boolean;
  signal next_add_dest_dim0_734_592_buf_req_0 : boolean;
  signal next_add_dest_dim0_734_592_buf_ack_0 : boolean;
  signal next_add_dest_dim0_734_592_buf_req_1 : boolean;
  signal next_add_dest_dim0_734_592_buf_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_875_inst_ack_0 : boolean;
  signal phi_stmt_593_req_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal phi_stmt_593_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_875_inst_req_0 : boolean;
  signal array_obj_ref_956_index_offset_ack_1 : boolean;
  signal phi_stmt_593_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_872_inst_ack_1 : boolean;
  signal add_dest_dim1_init_570_595_buf_req_0 : boolean;
  signal add_dest_dim1_init_570_595_buf_ack_0 : boolean;
  signal type_cast_807_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_872_inst_req_1 : boolean;
  signal add_dest_dim1_init_570_595_buf_req_1 : boolean;
  signal add_dest_dim1_init_570_595_buf_ack_1 : boolean;
  signal next_add_dest_dim1_728_596_buf_req_0 : boolean;
  signal next_add_dest_dim1_728_596_buf_ack_0 : boolean;
  signal ptr_deref_961_load_0_ack_0 : boolean;
  signal next_add_dest_dim1_728_596_buf_req_1 : boolean;
  signal next_add_dest_dim1_728_596_buf_ack_1 : boolean;
  signal type_cast_807_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_872_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_872_inst_req_0 : boolean;
  signal phi_stmt_597_req_1 : boolean;
  signal phi_stmt_597_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_869_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_869_inst_req_1 : boolean;
  signal phi_stmt_597_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_869_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_869_inst_req_0 : boolean;
  signal type_cast_867_inst_ack_1 : boolean;
  signal type_cast_867_inst_req_1 : boolean;
  signal type_cast_867_inst_ack_0 : boolean;
  signal type_cast_867_inst_req_0 : boolean;
  signal next_add_src_715_600_buf_req_0 : boolean;
  signal next_add_src_715_600_buf_ack_0 : boolean;
  signal type_cast_807_inst_req_0 : boolean;
  signal next_add_src_715_600_buf_req_1 : boolean;
  signal next_add_src_715_600_buf_ack_1 : boolean;
  signal type_cast_857_inst_ack_1 : boolean;
  signal type_cast_857_inst_req_1 : boolean;
  signal type_cast_857_inst_ack_0 : boolean;
  signal type_cast_857_inst_req_0 : boolean;
  signal ptr_deref_961_load_0_ack_1 : boolean;
  signal type_cast_847_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_1 : boolean;
  signal ptr_deref_961_load_0_req_1 : boolean;
  signal call_stmt_777_call_ack_0 : boolean;
  signal array_obj_ref_632_index_offset_req_0 : boolean;
  signal if_stmt_900_branch_ack_0 : boolean;
  signal array_obj_ref_632_index_offset_ack_0 : boolean;
  signal array_obj_ref_632_index_offset_req_1 : boolean;
  signal array_obj_ref_632_index_offset_ack_1 : boolean;
  signal if_stmt_900_branch_ack_1 : boolean;
  signal addr_of_633_final_reg_req_0 : boolean;
  signal addr_of_633_final_reg_ack_0 : boolean;
  signal call_stmt_777_call_req_0 : boolean;
  signal addr_of_633_final_reg_req_1 : boolean;
  signal addr_of_633_final_reg_ack_1 : boolean;
  signal ptr_deref_637_load_0_req_0 : boolean;
  signal ptr_deref_637_load_0_ack_0 : boolean;
  signal ptr_deref_637_load_0_req_1 : boolean;
  signal ptr_deref_637_load_0_ack_1 : boolean;
  signal array_obj_ref_644_index_offset_req_0 : boolean;
  signal array_obj_ref_644_index_offset_ack_0 : boolean;
  signal array_obj_ref_644_index_offset_req_1 : boolean;
  signal array_obj_ref_644_index_offset_ack_1 : boolean;
  signal addr_of_645_final_reg_req_0 : boolean;
  signal addr_of_645_final_reg_ack_0 : boolean;
  signal addr_of_645_final_reg_req_1 : boolean;
  signal addr_of_645_final_reg_ack_1 : boolean;
  signal W_ov_647_delayed_6_0_647_inst_req_0 : boolean;
  signal W_ov_647_delayed_6_0_647_inst_ack_0 : boolean;
  signal W_ov_647_delayed_6_0_647_inst_req_1 : boolean;
  signal W_ov_647_delayed_6_0_647_inst_ack_1 : boolean;
  signal ptr_deref_651_store_0_req_0 : boolean;
  signal ptr_deref_651_store_0_ack_0 : boolean;
  signal ptr_deref_651_store_0_req_1 : boolean;
  signal ptr_deref_651_store_0_ack_1 : boolean;
  signal W_dim2_limit_658_delayed_1_0_659_inst_req_0 : boolean;
  signal W_dim2_limit_658_delayed_1_0_659_inst_ack_0 : boolean;
  signal W_dim2_limit_658_delayed_1_0_659_inst_req_1 : boolean;
  signal W_dim2_limit_658_delayed_1_0_659_inst_ack_1 : boolean;
  signal SUB_u16_u16_670_inst_req_0 : boolean;
  signal SUB_u16_u16_670_inst_ack_0 : boolean;
  signal SUB_u16_u16_670_inst_req_1 : boolean;
  signal SUB_u16_u16_670_inst_ack_1 : boolean;
  signal W_nid1_true4_711_delayed_1_0_716_inst_req_0 : boolean;
  signal W_nid1_true4_711_delayed_1_0_716_inst_ack_0 : boolean;
  signal W_nid1_true4_711_delayed_1_0_716_inst_req_1 : boolean;
  signal W_nid1_true4_711_delayed_1_0_716_inst_ack_1 : boolean;
  signal SUB_u16_u16_760_inst_req_0 : boolean;
  signal SUB_u16_u16_760_inst_ack_0 : boolean;
  signal SUB_u16_u16_760_inst_req_1 : boolean;
  signal SUB_u16_u16_760_inst_ack_1 : boolean;
  signal do_while_stmt_575_branch_ack_0 : boolean;
  signal do_while_stmt_575_branch_ack_1 : boolean;
  signal type_cast_965_inst_req_0 : boolean;
  signal type_cast_965_inst_ack_0 : boolean;
  signal type_cast_965_inst_req_1 : boolean;
  signal type_cast_965_inst_ack_1 : boolean;
  signal type_cast_975_inst_req_0 : boolean;
  signal type_cast_975_inst_ack_0 : boolean;
  signal type_cast_975_inst_req_1 : boolean;
  signal type_cast_975_inst_ack_1 : boolean;
  signal type_cast_985_inst_req_0 : boolean;
  signal type_cast_985_inst_ack_0 : boolean;
  signal type_cast_985_inst_req_1 : boolean;
  signal type_cast_985_inst_ack_1 : boolean;
  signal type_cast_995_inst_req_0 : boolean;
  signal type_cast_995_inst_ack_0 : boolean;
  signal type_cast_995_inst_req_1 : boolean;
  signal type_cast_995_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_0 : boolean;
  signal type_cast_1005_inst_ack_0 : boolean;
  signal type_cast_1005_inst_req_1 : boolean;
  signal type_cast_1005_inst_ack_1 : boolean;
  signal type_cast_1015_inst_req_0 : boolean;
  signal type_cast_1015_inst_ack_0 : boolean;
  signal type_cast_1015_inst_req_1 : boolean;
  signal type_cast_1015_inst_ack_1 : boolean;
  signal type_cast_1025_inst_req_0 : boolean;
  signal type_cast_1025_inst_ack_0 : boolean;
  signal type_cast_1025_inst_req_1 : boolean;
  signal type_cast_1025_inst_ack_1 : boolean;
  signal type_cast_1035_inst_req_0 : boolean;
  signal type_cast_1035_inst_ack_0 : boolean;
  signal type_cast_1035_inst_req_1 : boolean;
  signal type_cast_1035_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1037_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1037_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1037_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1037_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1040_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1040_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1040_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1040_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1043_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1043_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1043_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1043_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1046_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1046_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1046_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1046_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1049_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1049_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1049_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1049_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1052_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1052_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1052_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1052_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1055_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1055_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1055_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1055_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1058_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1058_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1058_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1058_inst_ack_1 : boolean;
  signal if_stmt_1072_branch_req_0 : boolean;
  signal if_stmt_1072_branch_ack_1 : boolean;
  signal if_stmt_1072_branch_ack_0 : boolean;
  signal phi_stmt_282_req_0 : boolean;
  signal type_cast_288_inst_req_0 : boolean;
  signal type_cast_288_inst_ack_0 : boolean;
  signal type_cast_288_inst_req_1 : boolean;
  signal type_cast_288_inst_ack_1 : boolean;
  signal phi_stmt_282_req_1 : boolean;
  signal phi_stmt_282_ack_0 : boolean;
  signal phi_stmt_502_req_0 : boolean;
  signal type_cast_508_inst_req_0 : boolean;
  signal type_cast_508_inst_ack_0 : boolean;
  signal type_cast_508_inst_req_1 : boolean;
  signal type_cast_508_inst_ack_1 : boolean;
  signal phi_stmt_502_req_1 : boolean;
  signal phi_stmt_502_ack_0 : boolean;
  signal phi_stmt_944_req_0 : boolean;
  signal type_cast_950_inst_req_0 : boolean;
  signal type_cast_950_inst_ack_0 : boolean;
  signal type_cast_950_inst_req_1 : boolean;
  signal type_cast_950_inst_ack_1 : boolean;
  signal phi_stmt_944_req_1 : boolean;
  signal phi_stmt_944_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad_same_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad_same_CP_159_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad_same_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_same_CP_159_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad_same_CP_159_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_same_CP_159_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad_same_CP_159: Block -- control-path 
    signal zeropad_same_CP_159_elements: BooleanArray(415 downto 0);
    -- 
  begin -- 
    zeropad_same_CP_159_elements(0) <= zeropad_same_CP_159_start;
    zeropad_same_CP_159_symbol <= zeropad_same_CP_159_elements(415);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	29 
    -- CP-element group 0:  members (56) 
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_38/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/branch_block_stmt_38__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Update/cr
      -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_58_inst_req_1); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_0); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_45_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_70_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_83_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_95_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_108_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_120_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_133_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_145_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_158_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_170_inst_req_1); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_183_inst_req_1); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_193_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_202_inst_req_1); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(0), ack => type_cast_220_inst_req_1); -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	296 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	297 
    -- CP-element group 1: 	298 
    -- CP-element group 1: 	299 
    -- CP-element group 1: 	300 
    -- CP-element group 1: 	302 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_38/do_while_stmt_575__exit__
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793__entry__
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_update_start_
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_update_start_
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Update/ccr
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Sample/crr
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_update_start_
      -- CP-element group 1: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Sample/$entry
      -- 
    cr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(1), ack => type_cast_787_inst_req_1); -- 
    ccr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(1), ack => call_stmt_777_call_req_1); -- 
    cr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(1), ack => type_cast_782_inst_req_1); -- 
    rr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(1), ack => type_cast_782_inst_req_0); -- 
    crr_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(1), ack => call_stmt_777_call_req_0); -- 
    zeropad_same_CP_159_elements(1) <= zeropad_same_CP_159_elements(296);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_update_start_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_0, ack => zeropad_same_CP_159_elements(2)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(2), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_40_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_1, ack => zeropad_same_CP_159_elements(3)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(3), ack => type_cast_45_inst_req_0); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(3), ack => RPIPE_ConvTranspose_input_pipe_54_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_0, ack => zeropad_same_CP_159_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	53 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_45_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_1, ack => zeropad_same_CP_159_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_update_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_54_inst_ack_0, ack => zeropad_same_CP_159_elements(6)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(6), ack => RPIPE_ConvTranspose_input_pipe_54_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_54_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_54_inst_ack_1, ack => zeropad_same_CP_159_elements(7)); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(7), ack => type_cast_58_inst_req_0); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(7), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_0, ack => zeropad_same_CP_159_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	53 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_58_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_1, ack => zeropad_same_CP_159_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_update_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_0, ack => zeropad_same_CP_159_elements(10)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(10), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_66_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_1, ack => zeropad_same_CP_159_elements(11)); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(11), ack => type_cast_70_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(11), ack => RPIPE_ConvTranspose_input_pipe_79_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_0, ack => zeropad_same_CP_159_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	53 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_70_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_1, ack => zeropad_same_CP_159_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_update_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_79_inst_ack_0, ack => zeropad_same_CP_159_elements(14)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(14), ack => RPIPE_ConvTranspose_input_pipe_79_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_79_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Sample/rr
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_79_inst_ack_1, ack => zeropad_same_CP_159_elements(15)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(15), ack => type_cast_83_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(15), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => zeropad_same_CP_159_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	53 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_83_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => zeropad_same_CP_159_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_update_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Update/cr
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_0, ack => zeropad_same_CP_159_elements(18)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(18), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_91_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_1, ack => zeropad_same_CP_159_elements(19)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(19), ack => type_cast_95_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(19), ack => RPIPE_ConvTranspose_input_pipe_104_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => zeropad_same_CP_159_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	50 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_95_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => zeropad_same_CP_159_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_update_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_104_inst_ack_0, ack => zeropad_same_CP_159_elements(22)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(22), ack => RPIPE_ConvTranspose_input_pipe_104_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_104_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_104_inst_ack_1, ack => zeropad_same_CP_159_elements(23)); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(23), ack => type_cast_108_inst_req_0); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(23), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_0, ack => zeropad_same_CP_159_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25: 	56 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_108_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_1, ack => zeropad_same_CP_159_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_update_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_0, ack => zeropad_same_CP_159_elements(26)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(26), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_116_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_1, ack => zeropad_same_CP_159_elements(27)); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(27), ack => type_cast_120_inst_req_0); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(27), ack => RPIPE_ConvTranspose_input_pipe_129_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_0, ack => zeropad_same_CP_159_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	59 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_120_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_1, ack => zeropad_same_CP_159_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_update_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_129_inst_ack_0, ack => zeropad_same_CP_159_elements(30)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(30), ack => RPIPE_ConvTranspose_input_pipe_129_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_129_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_129_inst_ack_1, ack => zeropad_same_CP_159_elements(31)); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(31), ack => type_cast_133_inst_req_0); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(31), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_133_inst_ack_0, ack => zeropad_same_CP_159_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	59 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_133_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_133_inst_ack_1, ack => zeropad_same_CP_159_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_update_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_0, ack => zeropad_same_CP_159_elements(34)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(34), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_141_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_1, ack => zeropad_same_CP_159_elements(35)); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(35), ack => RPIPE_ConvTranspose_input_pipe_154_inst_req_0); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(35), ack => type_cast_145_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_0, ack => zeropad_same_CP_159_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	59 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_145_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_1, ack => zeropad_same_CP_159_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_update_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_154_inst_ack_0, ack => zeropad_same_CP_159_elements(38)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(38), ack => RPIPE_ConvTranspose_input_pipe_154_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_154_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_154_inst_ack_1, ack => zeropad_same_CP_159_elements(39)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(39), ack => type_cast_158_inst_req_0); -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(39), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_158_inst_ack_0, ack => zeropad_same_CP_159_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	59 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_158_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_158_inst_ack_1, ack => zeropad_same_CP_159_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_update_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Update/cr
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_0, ack => zeropad_same_CP_159_elements(42)); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(42), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_166_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Sample/rr
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_1, ack => zeropad_same_CP_159_elements(43)); -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(43), ack => RPIPE_ConvTranspose_input_pipe_179_inst_req_0); -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(43), ack => type_cast_170_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_0, ack => zeropad_same_CP_159_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	62 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_170_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_1, ack => zeropad_same_CP_159_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_update_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Update/cr
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_179_inst_ack_0, ack => zeropad_same_CP_159_elements(46)); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(46), ack => RPIPE_ConvTranspose_input_pipe_179_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/RPIPE_ConvTranspose_input_pipe_179_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Sample/rr
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_179_inst_ack_1, ack => zeropad_same_CP_159_elements(47)); -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(47), ack => type_cast_183_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Sample/ra
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_183_inst_ack_0, ack => zeropad_same_CP_159_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	62 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_183_Update/ca
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_183_inst_ack_1, ack => zeropad_same_CP_159_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	21 
    -- CP-element group 50: 	25 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Sample/rr
      -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(50), ack => type_cast_193_inst_req_0); -- 
    zeropad_same_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(21) & zeropad_same_CP_159_elements(25);
      gj_zeropad_same_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Sample/ra
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_0, ack => zeropad_same_CP_159_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	62 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_193_Update/ca
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_1, ack => zeropad_same_CP_159_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	5 
    -- CP-element group 53: 	9 
    -- CP-element group 53: 	13 
    -- CP-element group 53: 	17 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Sample/rr
      -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(53), ack => type_cast_202_inst_req_0); -- 
    zeropad_same_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(5) & zeropad_same_CP_159_elements(9) & zeropad_same_CP_159_elements(13) & zeropad_same_CP_159_elements(17);
      gj_zeropad_same_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_0, ack => zeropad_same_CP_159_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	62 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_202_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_1, ack => zeropad_same_CP_159_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	25 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Sample/rr
      -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(56), ack => type_cast_211_inst_req_0); -- 
    zeropad_same_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(21) & zeropad_same_CP_159_elements(25);
      gj_zeropad_same_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Sample/ra
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => zeropad_same_CP_159_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	62 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_211_Update/ca
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => zeropad_same_CP_159_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	33 
    -- CP-element group 59: 	41 
    -- CP-element group 59: 	37 
    -- CP-element group 59: 	29 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Sample/rr
      -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(59), ack => type_cast_220_inst_req_0); -- 
    zeropad_same_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(33) & zeropad_same_CP_159_elements(41) & zeropad_same_CP_159_elements(37) & zeropad_same_CP_159_elements(29);
      gj_zeropad_same_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Sample/ra
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_0, ack => zeropad_same_CP_159_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/type_cast_220_Update/ca
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_1, ack => zeropad_same_CP_159_elements(61)); -- 
    -- CP-element group 62:  branch  join  transition  place  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	49 
    -- CP-element group 62: 	45 
    -- CP-element group 62: 	52 
    -- CP-element group 62: 	61 
    -- CP-element group 62: 	55 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (10) 
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233__exit__
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234__entry__
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_233/$exit
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_38/R_cmp467_235_place
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_38/if_stmt_234_else_link/$entry
      -- 
    branch_req_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(62), ack => if_stmt_234_branch_req_0); -- 
    zeropad_same_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(49) & zeropad_same_CP_159_elements(45) & zeropad_same_CP_159_elements(52) & zeropad_same_CP_159_elements(61) & zeropad_same_CP_159_elements(55) & zeropad_same_CP_159_elements(58);
      gj_zeropad_same_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 branch_block_stmt_38/merge_stmt_244__exit__
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279__entry__
      -- CP-element group 63: 	 branch_block_stmt_38/if_stmt_234_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_38/if_stmt_234_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_38/entry_bbx_xnph469
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_update_start_
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_38/entry_bbx_xnph469_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/entry_bbx_xnph469_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_38/merge_stmt_244_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_38/merge_stmt_244_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/merge_stmt_244_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_38/merge_stmt_244_PhiAck/dummy
      -- 
    if_choice_transition_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_234_branch_ack_1, ack => zeropad_same_CP_159_elements(63)); -- 
    rr_659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(63), ack => type_cast_265_inst_req_0); -- 
    cr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(63), ack => type_cast_265_inst_req_1); -- 
    -- CP-element group 64:  transition  place  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	395 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_38/if_stmt_234_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_38/if_stmt_234_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_38/entry_forx_xcond171x_xpreheader
      -- CP-element group 64: 	 branch_block_stmt_38/entry_forx_xcond171x_xpreheader_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_38/entry_forx_xcond171x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_234_branch_ack_0, ack => zeropad_same_CP_159_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Sample/ra
      -- 
    ra_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_0, ack => zeropad_same_CP_159_elements(65)); -- 
    -- CP-element group 66:  transition  place  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	396 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279__exit__
      -- CP-element group 66: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/$exit
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_250_to_assign_stmt_279/type_cast_265_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_282/$entry
      -- CP-element group 66: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/$entry
      -- 
    ca_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_1, ack => zeropad_same_CP_159_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	401 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	106 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Sample/ack
      -- 
    ack_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_294_index_offset_ack_0, ack => zeropad_same_CP_159_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	401 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_request/req
      -- 
    ack_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_294_index_offset_ack_1, ack => zeropad_same_CP_159_elements(68)); -- 
    req_708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(68), ack => addr_of_295_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_request/ack
      -- 
    ack_709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_295_final_reg_ack_0, ack => zeropad_same_CP_159_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	401 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	103 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_word_addrgen/root_register_ack
      -- 
    ack_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_295_final_reg_ack_1, ack => zeropad_same_CP_159_elements(70)); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	401 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_update_start_
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Update/cr
      -- 
    ra_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_0, ack => zeropad_same_CP_159_elements(71)); -- 
    cr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(71), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (9) 
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Sample/rr
      -- 
    ca_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_1, ack => zeropad_same_CP_159_elements(72)); -- 
    rr_736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(72), ack => type_cast_302_inst_req_0); -- 
    rr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(72), ack => RPIPE_ConvTranspose_input_pipe_311_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Sample/ra
      -- 
    ra_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_0, ack => zeropad_same_CP_159_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	401 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	103 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Update/ca
      -- 
    ca_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_1, ack => zeropad_same_CP_159_elements(74)); -- 
    -- CP-element group 75:  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (6) 
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_update_start_
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Update/cr
      -- 
    ra_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_311_inst_ack_0, ack => zeropad_same_CP_159_elements(75)); -- 
    cr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(75), ack => RPIPE_ConvTranspose_input_pipe_311_inst_req_1); -- 
    -- CP-element group 76:  fork  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	79 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_311_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Sample/rr
      -- 
    ca_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_311_inst_ack_1, ack => zeropad_same_CP_159_elements(76)); -- 
    rr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(76), ack => type_cast_315_inst_req_0); -- 
    rr_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(76), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_0); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Sample/ra
      -- 
    ra_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_0, ack => zeropad_same_CP_159_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	401 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	103 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Update/ca
      -- 
    ca_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_1, ack => zeropad_same_CP_159_elements(78)); -- 
    -- CP-element group 79:  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	76 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_update_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Update/cr
      -- 
    ra_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_0, ack => zeropad_same_CP_159_elements(79)); -- 
    cr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(79), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_329_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Sample/rr
      -- 
    ca_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_1, ack => zeropad_same_CP_159_elements(80)); -- 
    rr_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(80), ack => type_cast_333_inst_req_0); -- 
    rr_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(80), ack => RPIPE_ConvTranspose_input_pipe_347_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Sample/ra
      -- 
    ra_793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_0, ack => zeropad_same_CP_159_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	401 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	103 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Update/ca
      -- 
    ca_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_1, ack => zeropad_same_CP_159_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_update_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Update/cr
      -- 
    ra_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_347_inst_ack_0, ack => zeropad_same_CP_159_elements(83)); -- 
    cr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(83), ack => RPIPE_ConvTranspose_input_pipe_347_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	87 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_347_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Sample/rr
      -- 
    ca_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_347_inst_ack_1, ack => zeropad_same_CP_159_elements(84)); -- 
    rr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(84), ack => type_cast_351_inst_req_0); -- 
    rr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(84), ack => RPIPE_ConvTranspose_input_pipe_365_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Sample/ra
      -- 
    ra_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_351_inst_ack_0, ack => zeropad_same_CP_159_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	401 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	103 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Update/ca
      -- 
    ca_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_351_inst_ack_1, ack => zeropad_same_CP_159_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	84 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_update_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Update/cr
      -- 
    ra_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_365_inst_ack_0, ack => zeropad_same_CP_159_elements(87)); -- 
    cr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(87), ack => RPIPE_ConvTranspose_input_pipe_365_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	91 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_365_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Sample/rr
      -- 
    ca_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_365_inst_ack_1, ack => zeropad_same_CP_159_elements(88)); -- 
    rr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(88), ack => type_cast_369_inst_req_0); -- 
    rr_862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(88), ack => RPIPE_ConvTranspose_input_pipe_383_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Sample/ra
      -- 
    ra_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_369_inst_ack_0, ack => zeropad_same_CP_159_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	401 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	103 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Update/ca
      -- 
    ca_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_369_inst_ack_1, ack => zeropad_same_CP_159_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_update_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Update/cr
      -- 
    ra_863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_383_inst_ack_0, ack => zeropad_same_CP_159_elements(91)); -- 
    cr_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(91), ack => RPIPE_ConvTranspose_input_pipe_383_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_383_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Sample/rr
      -- 
    ca_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_383_inst_ack_1, ack => zeropad_same_CP_159_elements(92)); -- 
    rr_876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(92), ack => type_cast_387_inst_req_0); -- 
    rr_890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(92), ack => RPIPE_ConvTranspose_input_pipe_401_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Sample/ra
      -- 
    ra_877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_387_inst_ack_0, ack => zeropad_same_CP_159_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	401 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	103 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Update/ca
      -- 
    ca_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_387_inst_ack_1, ack => zeropad_same_CP_159_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_update_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Update/cr
      -- 
    ra_891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_401_inst_ack_0, ack => zeropad_same_CP_159_elements(95)); -- 
    cr_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(95), ack => RPIPE_ConvTranspose_input_pipe_401_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_401_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Sample/rr
      -- 
    ca_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_401_inst_ack_1, ack => zeropad_same_CP_159_elements(96)); -- 
    rr_904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(96), ack => type_cast_405_inst_req_0); -- 
    rr_918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(96), ack => RPIPE_ConvTranspose_input_pipe_419_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Sample/ra
      -- 
    ra_905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_405_inst_ack_0, ack => zeropad_same_CP_159_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	401 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Update/ca
      -- 
    ca_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_405_inst_ack_1, ack => zeropad_same_CP_159_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_update_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Update/cr
      -- 
    ra_919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_419_inst_ack_0, ack => zeropad_same_CP_159_elements(99)); -- 
    cr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(99), ack => RPIPE_ConvTranspose_input_pipe_419_inst_req_1); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_419_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Sample/rr
      -- 
    ca_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_419_inst_ack_1, ack => zeropad_same_CP_159_elements(100)); -- 
    rr_932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(100), ack => type_cast_423_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Sample/ra
      -- 
    ra_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_423_inst_ack_0, ack => zeropad_same_CP_159_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	401 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Update/ca
      -- 
    ca_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_423_inst_ack_1, ack => zeropad_same_CP_159_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	70 
    -- CP-element group 103: 	74 
    -- CP-element group 103: 	78 
    -- CP-element group 103: 	82 
    -- CP-element group 103: 	86 
    -- CP-element group 103: 	90 
    -- CP-element group 103: 	94 
    -- CP-element group 103: 	98 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/ptr_deref_431_Split/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/ptr_deref_431_Split/$exit
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/ptr_deref_431_Split/split_req
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/ptr_deref_431_Split/split_ack
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/word_access_start/word_0/rr
      -- 
    rr_976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(103), ack => ptr_deref_431_store_0_req_0); -- 
    zeropad_same_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(70) & zeropad_same_CP_159_elements(74) & zeropad_same_CP_159_elements(78) & zeropad_same_CP_159_elements(82) & zeropad_same_CP_159_elements(86) & zeropad_same_CP_159_elements(90) & zeropad_same_CP_159_elements(94) & zeropad_same_CP_159_elements(98) & zeropad_same_CP_159_elements(102);
      gj_zeropad_same_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/word_access_start/$exit
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/word_access_start/word_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Sample/word_access_start/word_0/ra
      -- 
    ra_977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_431_store_0_ack_0, ack => zeropad_same_CP_159_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	401 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/word_access_complete/$exit
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/word_access_complete/word_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/word_access_complete/word_0/ca
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_431_store_0_ack_1, ack => zeropad_same_CP_159_elements(105)); -- 
    -- CP-element group 106:  branch  join  transition  place  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	67 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (10) 
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444__exit__
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445__entry__
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/$exit
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445_dead_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445_eval_test/$entry
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445_eval_test/$exit
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445_eval_test/branch_req
      -- CP-element group 106: 	 branch_block_stmt_38/R_exitcond2_446_place
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445_if_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_38/if_stmt_445_else_link/$entry
      -- 
    branch_req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(106), ack => if_stmt_445_branch_req_0); -- 
    zeropad_same_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(67) & zeropad_same_CP_159_elements(105);
      gj_zeropad_same_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  merge  transition  place  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	395 
    -- CP-element group 107:  members (13) 
      -- CP-element group 107: 	 branch_block_stmt_38/merge_stmt_240__exit__
      -- CP-element group 107: 	 branch_block_stmt_38/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader
      -- CP-element group 107: 	 branch_block_stmt_38/if_stmt_445_if_link/$exit
      -- CP-element group 107: 	 branch_block_stmt_38/if_stmt_445_if_link/if_choice_transition
      -- CP-element group 107: 	 branch_block_stmt_38/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit
      -- CP-element group 107: 	 branch_block_stmt_38/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 107: 	 branch_block_stmt_38/merge_stmt_240_PhiReqMerge
      -- CP-element group 107: 	 branch_block_stmt_38/merge_stmt_240_PhiAck/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/merge_stmt_240_PhiAck/$exit
      -- CP-element group 107: 	 branch_block_stmt_38/merge_stmt_240_PhiAck/dummy
      -- CP-element group 107: 	 branch_block_stmt_38/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_445_branch_ack_1, ack => zeropad_same_CP_159_elements(107)); -- 
    -- CP-element group 108:  fork  transition  place  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	397 
    -- CP-element group 108: 	398 
    -- CP-element group 108:  members (12) 
      -- CP-element group 108: 	 branch_block_stmt_38/if_stmt_445_else_link/$exit
      -- CP-element group 108: 	 branch_block_stmt_38/if_stmt_445_else_link/else_choice_transition
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_445_branch_ack_0, ack => zeropad_same_CP_159_elements(108)); -- 
    rr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(108), ack => type_cast_288_inst_req_0); -- 
    cr_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(108), ack => type_cast_288_inst_req_1); -- 
    -- CP-element group 109:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	395 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (18) 
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_update_start_
      -- CP-element group 109: 	 branch_block_stmt_38/merge_stmt_464__exit__
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499__entry__
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/$entry
      -- CP-element group 109: 	 branch_block_stmt_38/if_stmt_458_if_link/if_choice_transition
      -- CP-element group 109: 	 branch_block_stmt_38/forx_xend250_bbx_xnph450
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_38/if_stmt_458_if_link/$exit
      -- CP-element group 109: 	 branch_block_stmt_38/forx_xend250_bbx_xnph450_PhiReq/$entry
      -- CP-element group 109: 	 branch_block_stmt_38/forx_xend250_bbx_xnph450_PhiReq/$exit
      -- CP-element group 109: 	 branch_block_stmt_38/merge_stmt_464_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_38/merge_stmt_464_PhiAck/$entry
      -- CP-element group 109: 	 branch_block_stmt_38/merge_stmt_464_PhiAck/$exit
      -- CP-element group 109: 	 branch_block_stmt_38/merge_stmt_464_PhiAck/dummy
      -- 
    if_choice_transition_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_458_branch_ack_1, ack => zeropad_same_CP_159_elements(109)); -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(109), ack => type_cast_485_inst_req_1); -- 
    rr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(109), ack => type_cast_485_inst_req_0); -- 
    -- CP-element group 110:  transition  place  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	395 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	408 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_38/forx_xend250_forx_xend273
      -- CP-element group 110: 	 branch_block_stmt_38/if_stmt_458_else_link/else_choice_transition
      -- CP-element group 110: 	 branch_block_stmt_38/if_stmt_458_else_link/$exit
      -- CP-element group 110: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 110: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_458_branch_ack_0, ack => zeropad_same_CP_159_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Sample/ra
      -- 
    ra_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_0, ack => zeropad_same_CP_159_elements(111)); -- 
    -- CP-element group 112:  transition  place  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	402 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499__exit__
      -- CP-element group 112: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/$exit
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_470_to_assign_stmt_499/type_cast_485_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/$entry
      -- CP-element group 112: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_502/$entry
      -- CP-element group 112: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/$entry
      -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_1, ack => zeropad_same_CP_159_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	407 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	119 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_sample_complete
      -- 
    ack_1075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_514_index_offset_ack_0, ack => zeropad_same_CP_159_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	407 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (11) 
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_base_plus_offset/sum_rename_ack
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_request/req
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_request/$entry
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_base_plus_offset/sum_rename_req
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_base_plus_offset/$exit
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_base_plus_offset/$entry
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Update/ack
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_offset_calculated
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_root_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_sample_start_
      -- 
    ack_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_514_index_offset_ack_1, ack => zeropad_same_CP_159_elements(114)); -- 
    req_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(114), ack => addr_of_515_final_reg_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_request/ack
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_request/$exit
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_sample_completed_
      -- 
    ack_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_515_final_reg_ack_0, ack => zeropad_same_CP_159_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	407 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (28) 
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_plus_offset/sum_rename_req
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_plus_offset/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_complete/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_plus_offset/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_addr_resize/base_resize_ack
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_addr_resize/base_resize_req
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_addr_resize/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_addr_resize/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_address_resized
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_complete/ack
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/ptr_deref_518_Split/split_ack
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/ptr_deref_518_Split/split_req
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/ptr_deref_518_Split/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/ptr_deref_518_Split/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_word_addrgen/root_register_ack
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_word_addrgen/root_register_req
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_word_addrgen/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_word_addrgen/$entry
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_base_plus_offset/sum_rename_ack
      -- 
    ack_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_515_final_reg_ack_1, ack => zeropad_same_CP_159_elements(116)); -- 
    rr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(116), ack => ptr_deref_518_store_0_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/word_access_start/word_0/ra
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Sample/$exit
      -- 
    ra_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_518_store_0_ack_0, ack => zeropad_same_CP_159_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	407 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/$exit
      -- 
    ca_1145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_518_store_0_ack_1, ack => zeropad_same_CP_159_elements(118)); -- 
    -- CP-element group 119:  branch  join  transition  place  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	113 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (10) 
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533_if_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533_eval_test/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533_eval_test/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533_dead_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/R_exitcond_534_place
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532__exit__
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533__entry__
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533_eval_test/branch_req
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_533_else_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/$exit
      -- 
    branch_req_1153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(119), ack => if_stmt_533_branch_req_0); -- 
    zeropad_same_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(113) & zeropad_same_CP_159_elements(118);
      gj_zeropad_same_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  merge  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	408 
    -- CP-element group 120:  members (13) 
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_533_if_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_38/merge_stmt_539__exit__
      -- CP-element group 120: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 120: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_533_if_link/if_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 120: 	 branch_block_stmt_38/merge_stmt_539_PhiReqMerge
      -- CP-element group 120: 	 branch_block_stmt_38/merge_stmt_539_PhiAck/$entry
      -- CP-element group 120: 	 branch_block_stmt_38/merge_stmt_539_PhiAck/$exit
      -- CP-element group 120: 	 branch_block_stmt_38/merge_stmt_539_PhiAck/dummy
      -- CP-element group 120: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_533_branch_ack_1, ack => zeropad_same_CP_159_elements(120)); -- 
    -- CP-element group 121:  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	403 
    -- CP-element group 121: 	404 
    -- CP-element group 121:  members (12) 
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_533_else_link/else_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_533_else_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_533_branch_ack_0, ack => zeropad_same_CP_159_elements(121)); -- 
    rr_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(121), ack => type_cast_508_inst_req_0); -- 
    cr_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(121), ack => type_cast_508_inst_req_1); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	408 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Sample/cra
      -- CP-element group 122: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_sample_completed_
      -- 
    cra_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_544_call_ack_0, ack => zeropad_same_CP_159_elements(122)); -- 
    -- CP-element group 123:  transition  place  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	408 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (10) 
      -- CP-element group 123: 	 branch_block_stmt_38/call_stmt_544__exit__
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_549_to_assign_stmt_574__entry__
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_549_to_assign_stmt_574__exit__
      -- CP-element group 123: 	 branch_block_stmt_38/do_while_stmt_575__entry__
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_549_to_assign_stmt_574/$exit
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_549_to_assign_stmt_574/$entry
      -- CP-element group 123: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Update/cca
      -- CP-element group 123: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_38/call_stmt_544/$exit
      -- 
    cca_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_544_call_ack_1, ack => zeropad_same_CP_159_elements(123)); -- 
    -- CP-element group 124:  transition  place  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	130 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575__entry__
      -- CP-element group 124: 	 branch_block_stmt_38/do_while_stmt_575/$entry
      -- 
    zeropad_same_CP_159_elements(124) <= zeropad_same_CP_159_elements(123);
    -- CP-element group 125:  merge  place  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	296 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575__exit__
      -- 
    -- Element group zeropad_same_CP_159_elements(125) is bound as output of CP function.
    -- CP-element group 126:  merge  place  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	129 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_38/do_while_stmt_575/loop_back
      -- 
    -- Element group zeropad_same_CP_159_elements(126) is bound as output of CP function.
    -- CP-element group 127:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	132 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	294 
    -- CP-element group 127: 	295 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_38/do_while_stmt_575/condition_done
      -- CP-element group 127: 	 branch_block_stmt_38/do_while_stmt_575/loop_exit/$entry
      -- CP-element group 127: 	 branch_block_stmt_38/do_while_stmt_575/loop_taken/$entry
      -- 
    zeropad_same_CP_159_elements(127) <= zeropad_same_CP_159_elements(132);
    -- CP-element group 128:  branch  place  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	293 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_38/do_while_stmt_575/loop_body_done
      -- 
    zeropad_same_CP_159_elements(128) <= zeropad_same_CP_159_elements(293);
    -- CP-element group 129:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	141 
    -- CP-element group 129: 	160 
    -- CP-element group 129: 	179 
    -- CP-element group 129: 	198 
    -- CP-element group 129: 	217 
    -- CP-element group 129: 	236 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/back_edge_to_loop_body
      -- 
    zeropad_same_CP_159_elements(129) <= zeropad_same_CP_159_elements(126);
    -- CP-element group 130:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	124 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	143 
    -- CP-element group 130: 	162 
    -- CP-element group 130: 	181 
    -- CP-element group 130: 	200 
    -- CP-element group 130: 	219 
    -- CP-element group 130: 	238 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/first_time_through_loop_body
      -- 
    zeropad_same_CP_159_elements(130) <= zeropad_same_CP_159_elements(124);
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	137 
    -- CP-element group 131: 	138 
    -- CP-element group 131: 	154 
    -- CP-element group 131: 	155 
    -- CP-element group 131: 	173 
    -- CP-element group 131: 	174 
    -- CP-element group 131: 	192 
    -- CP-element group 131: 	193 
    -- CP-element group 131: 	211 
    -- CP-element group 131: 	212 
    -- CP-element group 131: 	230 
    -- CP-element group 131: 	231 
    -- CP-element group 131: 	250 
    -- CP-element group 131: 	251 
    -- CP-element group 131: 	261 
    -- CP-element group 131: 	263 
    -- CP-element group 131: 	276 
    -- CP-element group 131: 	280 
    -- CP-element group 131: 	284 
    -- CP-element group 131: 	288 
    -- CP-element group 131: 	292 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/loop_body_start
      -- CP-element group 131: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/$entry
      -- 
    -- Element group zeropad_same_CP_159_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	136 
    -- CP-element group 132: 	140 
    -- CP-element group 132: 	159 
    -- CP-element group 132: 	178 
    -- CP-element group 132: 	279 
    -- CP-element group 132: 	283 
    -- CP-element group 132: 	291 
    -- CP-element group 132: 	292 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	127 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/condition_evaluated
      -- 
    condition_evaluated_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(132), ack => do_while_stmt_575_branch_req_0); -- 
    zeropad_same_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(136) & zeropad_same_CP_159_elements(140) & zeropad_same_CP_159_elements(159) & zeropad_same_CP_159_elements(178) & zeropad_same_CP_159_elements(279) & zeropad_same_CP_159_elements(283) & zeropad_same_CP_159_elements(291) & zeropad_same_CP_159_elements(292);
      gj_zeropad_same_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	137 
    -- CP-element group 133: 	154 
    -- CP-element group 133: 	173 
    -- CP-element group 133: 	192 
    -- CP-element group 133: 	211 
    -- CP-element group 133: 	230 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	136 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	156 
    -- CP-element group 133: 	175 
    -- CP-element group 133: 	194 
    -- CP-element group 133: 	213 
    -- CP-element group 133: 	232 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/aggregated_phi_sample_req
      -- 
    zeropad_same_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(137) & zeropad_same_CP_159_elements(154) & zeropad_same_CP_159_elements(173) & zeropad_same_CP_159_elements(192) & zeropad_same_CP_159_elements(211) & zeropad_same_CP_159_elements(230) & zeropad_same_CP_159_elements(136);
      gj_zeropad_same_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	139 
    -- CP-element group 134: 	157 
    -- CP-element group 134: 	176 
    -- CP-element group 134: 	195 
    -- CP-element group 134: 	214 
    -- CP-element group 134: 	233 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	277 
    -- CP-element group 134: 	281 
    -- CP-element group 134: 	285 
    -- CP-element group 134: 	293 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134: 	154 
    -- CP-element group 134: 	173 
    -- CP-element group 134: 	192 
    -- CP-element group 134: 	211 
    -- CP-element group 134: 	230 
    -- CP-element group 134:  members (7) 
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/aggregated_phi_sample_ack
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_sample_completed_
      -- 
    zeropad_same_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(139) & zeropad_same_CP_159_elements(157) & zeropad_same_CP_159_elements(176) & zeropad_same_CP_159_elements(195) & zeropad_same_CP_159_elements(214) & zeropad_same_CP_159_elements(233);
      gj_zeropad_same_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	138 
    -- CP-element group 135: 	155 
    -- CP-element group 135: 	174 
    -- CP-element group 135: 	193 
    -- CP-element group 135: 	212 
    -- CP-element group 135: 	231 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	158 
    -- CP-element group 135: 	177 
    -- CP-element group 135: 	196 
    -- CP-element group 135: 	215 
    -- CP-element group 135: 	234 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/aggregated_phi_update_req
      -- CP-element group 135: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_update_start__ps
      -- 
    zeropad_same_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(138) & zeropad_same_CP_159_elements(155) & zeropad_same_CP_159_elements(174) & zeropad_same_CP_159_elements(193) & zeropad_same_CP_159_elements(212) & zeropad_same_CP_159_elements(231);
      gj_zeropad_same_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	140 
    -- CP-element group 136: 	159 
    -- CP-element group 136: 	178 
    -- CP-element group 136: 	197 
    -- CP-element group 136: 	216 
    -- CP-element group 136: 	235 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	132 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	133 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/aggregated_phi_update_ack
      -- 
    zeropad_same_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(140) & zeropad_same_CP_159_elements(159) & zeropad_same_CP_159_elements(178) & zeropad_same_CP_159_elements(197) & zeropad_same_CP_159_elements(216) & zeropad_same_CP_159_elements(235);
      gj_zeropad_same_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	131 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	279 
    -- CP-element group 137: 	283 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_sample_start_
      -- 
    zeropad_same_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(279) & zeropad_same_CP_159_elements(283);
      gj_zeropad_same_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	131 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	135 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_update_start_
      -- 
    zeropad_same_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(140);
      gj_zeropad_same_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	134 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	132 
    -- CP-element group 140: 	136 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_update_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	129 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_loopback_trigger
      -- 
    zeropad_same_CP_159_elements(141) <= zeropad_same_CP_159_elements(129);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_loopback_sample_req_ps
      -- CP-element group 142: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_loopback_sample_req
      -- 
    phi_stmt_577_loopback_sample_req_1214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_577_loopback_sample_req_1214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(142), ack => phi_stmt_577_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	130 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_entry_trigger
      -- 
    zeropad_same_CP_159_elements(143) <= zeropad_same_CP_159_elements(130);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_entry_sample_req_ps
      -- CP-element group 144: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_entry_sample_req
      -- 
    phi_stmt_577_entry_sample_req_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_577_entry_sample_req_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(144), ack => phi_stmt_577_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_phi_mux_ack_ps
      -- CP-element group 145: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_577_phi_mux_ack
      -- 
    phi_stmt_577_phi_mux_ack_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_577_ack_0, ack => zeropad_same_CP_159_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_sample_start__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_update_start_
      -- CP-element group 147: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_update_start__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_update_completed__ps
      -- 
    zeropad_same_CP_159_elements(148) <= zeropad_same_CP_159_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim0_init_579_update_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(147), ack => zeropad_same_CP_159_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_sample_start__ps
      -- 
    req_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(150), ack => next_input_dim0_756_580_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_update_start_
      -- CP-element group 151: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Update/req
      -- 
    req_1246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(151), ack => next_input_dim0_756_580_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_sample_completed__ps
      -- 
    ack_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_756_580_buf_ack_0, ack => zeropad_same_CP_159_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim0_580_Update/ack
      -- 
    ack_1247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_756_580_buf_ack_1, ack => zeropad_same_CP_159_elements(153)); -- 
    -- CP-element group 154:  join  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	131 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	134 
    -- CP-element group 154: 	279 
    -- CP-element group 154: 	283 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	133 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_sample_start_
      -- 
    zeropad_same_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(279) & zeropad_same_CP_159_elements(283);
      gj_zeropad_same_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	131 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	135 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_update_start_
      -- 
    zeropad_same_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(159);
      gj_zeropad_same_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	133 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_sample_start__ps
      -- 
    zeropad_same_CP_159_elements(156) <= zeropad_same_CP_159_elements(133);
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	134 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(157) is bound as output of CP function.
    -- CP-element group 158:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	135 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_update_start__ps
      -- 
    zeropad_same_CP_159_elements(158) <= zeropad_same_CP_159_elements(135);
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	132 
    -- CP-element group 159: 	136 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_update_completed__ps
      -- CP-element group 159: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_update_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(159) is bound as output of CP function.
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	129 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_loopback_trigger
      -- 
    zeropad_same_CP_159_elements(160) <= zeropad_same_CP_159_elements(129);
    -- CP-element group 161:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (2) 
      -- CP-element group 161: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_loopback_sample_req_ps
      -- CP-element group 161: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_loopback_sample_req
      -- 
    phi_stmt_581_loopback_sample_req_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_loopback_sample_req_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(161), ack => phi_stmt_581_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(161) is bound as output of CP function.
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	130 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_entry_trigger
      -- 
    zeropad_same_CP_159_elements(162) <= zeropad_same_CP_159_elements(130);
    -- CP-element group 163:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_entry_sample_req_ps
      -- CP-element group 163: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_entry_sample_req
      -- 
    phi_stmt_581_entry_sample_req_1261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_entry_sample_req_1261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(163), ack => phi_stmt_581_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(163) is bound as output of CP function.
    -- CP-element group 164:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_phi_mux_ack_ps
      -- CP-element group 164: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_581_phi_mux_ack
      -- 
    phi_stmt_581_phi_mux_ack_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_581_ack_0, ack => zeropad_same_CP_159_elements(164)); -- 
    -- CP-element group 165:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (4) 
      -- CP-element group 165: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_sample_completed__ps
      -- CP-element group 165: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_sample_start__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(165) is bound as output of CP function.
    -- CP-element group 166:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_update_start_
      -- CP-element group 166: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_update_start__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_update_completed__ps
      -- 
    zeropad_same_CP_159_elements(167) <= zeropad_same_CP_159_elements(168);
    -- CP-element group 168:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	167 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim1_init_583_update_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(168) is a control-delay.
    cp_element_168_delay: control_delay_element  generic map(name => " 168_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(166), ack => zeropad_same_CP_159_elements(168), clk => clk, reset =>reset);
    -- CP-element group 169:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (4) 
      -- CP-element group 169: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Sample/req
      -- CP-element group 169: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_sample_start__ps
      -- 
    req_1285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(169), ack => next_input_dim1_750_584_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Update/req
      -- CP-element group 170: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_update_start_
      -- CP-element group 170: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_update_start__ps
      -- 
    req_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(170), ack => next_input_dim1_750_584_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_sample_completed__ps
      -- 
    ack_1286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_750_584_buf_ack_0, ack => zeropad_same_CP_159_elements(171)); -- 
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim1_584_update_completed__ps
      -- 
    ack_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_750_584_buf_ack_1, ack => zeropad_same_CP_159_elements(172)); -- 
    -- CP-element group 173:  join  transition  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	131 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	134 
    -- CP-element group 173: 	279 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	133 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_sample_start_
      -- 
    zeropad_same_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(279);
      gj_zeropad_same_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	131 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	178 
    -- CP-element group 174: 	264 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	135 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_update_start_
      -- 
    zeropad_same_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(178) & zeropad_same_CP_159_elements(264);
      gj_zeropad_same_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	133 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_sample_start__ps
      -- 
    zeropad_same_CP_159_elements(175) <= zeropad_same_CP_159_elements(133);
    -- CP-element group 176:  join  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	134 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(176) is bound as output of CP function.
    -- CP-element group 177:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	135 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_update_start__ps
      -- 
    zeropad_same_CP_159_elements(177) <= zeropad_same_CP_159_elements(135);
    -- CP-element group 178:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	132 
    -- CP-element group 178: 	136 
    -- CP-element group 178: 	262 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	174 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_update_completed__ps
      -- CP-element group 178: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_update_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(178) is bound as output of CP function.
    -- CP-element group 179:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	129 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_loopback_trigger
      -- 
    zeropad_same_CP_159_elements(179) <= zeropad_same_CP_159_elements(129);
    -- CP-element group 180:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_loopback_sample_req_ps
      -- CP-element group 180: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_loopback_sample_req
      -- 
    phi_stmt_585_loopback_sample_req_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_loopback_sample_req_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(180), ack => phi_stmt_585_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(180) is bound as output of CP function.
    -- CP-element group 181:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	130 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_entry_trigger
      -- 
    zeropad_same_CP_159_elements(181) <= zeropad_same_CP_159_elements(130);
    -- CP-element group 182:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_entry_sample_req_ps
      -- CP-element group 182: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_entry_sample_req
      -- 
    phi_stmt_585_entry_sample_req_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_entry_sample_req_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(182), ack => phi_stmt_585_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(182) is bound as output of CP function.
    -- CP-element group 183:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_phi_mux_ack
      -- CP-element group 183: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_585_phi_mux_ack_ps
      -- 
    phi_stmt_585_phi_mux_ack_1308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_585_ack_0, ack => zeropad_same_CP_159_elements(183)); -- 
    -- CP-element group 184:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (4) 
      -- CP-element group 184: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_sample_completed__ps
      -- CP-element group 184: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_sample_start__ps
      -- CP-element group 184: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_sample_start_
      -- 
    -- Element group zeropad_same_CP_159_elements(184) is bound as output of CP function.
    -- CP-element group 185:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (2) 
      -- CP-element group 185: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_update_start__ps
      -- CP-element group 185: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_update_start_
      -- 
    -- Element group zeropad_same_CP_159_elements(185) is bound as output of CP function.
    -- CP-element group 186:  join  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_update_completed__ps
      -- 
    zeropad_same_CP_159_elements(186) <= zeropad_same_CP_159_elements(187);
    -- CP-element group 187:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	186 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_input_dim2_init_587_update_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(187) is a control-delay.
    cp_element_187_delay: control_delay_element  generic map(name => " 187_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(185), ack => zeropad_same_CP_159_elements(187), clk => clk, reset =>reset);
    -- CP-element group 188:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (4) 
      -- CP-element group 188: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Sample/req
      -- CP-element group 188: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_sample_start__ps
      -- 
    req_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(188), ack => next_input_dim2_740_588_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(188) is bound as output of CP function.
    -- CP-element group 189:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (4) 
      -- CP-element group 189: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_update_start__ps
      -- CP-element group 189: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Update/req
      -- CP-element group 189: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_update_start_
      -- CP-element group 189: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Update/$entry
      -- 
    req_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(189), ack => next_input_dim2_740_588_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(189) is bound as output of CP function.
    -- CP-element group 190:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (4) 
      -- CP-element group 190: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Sample/ack
      -- CP-element group 190: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_sample_completed__ps
      -- CP-element group 190: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Sample/$exit
      -- 
    ack_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_740_588_buf_ack_0, ack => zeropad_same_CP_159_elements(190)); -- 
    -- CP-element group 191:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (4) 
      -- CP-element group 191: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_update_completed__ps
      -- CP-element group 191: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Update/ack
      -- CP-element group 191: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_input_dim2_588_Update/$exit
      -- 
    ack_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_740_588_buf_ack_1, ack => zeropad_same_CP_159_elements(191)); -- 
    -- CP-element group 192:  join  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	131 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	134 
    -- CP-element group 192: 	279 
    -- CP-element group 192: 	283 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	133 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_sample_start_
      -- 
    zeropad_same_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(279) & zeropad_same_CP_159_elements(283);
      gj_zeropad_same_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	131 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	197 
    -- CP-element group 193: 	264 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	135 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_update_start_
      -- 
    zeropad_same_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(197) & zeropad_same_CP_159_elements(264);
      gj_zeropad_same_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	133 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_sample_start__ps
      -- 
    zeropad_same_CP_159_elements(194) <= zeropad_same_CP_159_elements(133);
    -- CP-element group 195:  join  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	134 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(195) is bound as output of CP function.
    -- CP-element group 196:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	135 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_update_start__ps
      -- 
    zeropad_same_CP_159_elements(196) <= zeropad_same_CP_159_elements(135);
    -- CP-element group 197:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	136 
    -- CP-element group 197: 	262 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	193 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_update_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(197) is bound as output of CP function.
    -- CP-element group 198:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	129 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_loopback_trigger
      -- 
    zeropad_same_CP_159_elements(198) <= zeropad_same_CP_159_elements(129);
    -- CP-element group 199:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_loopback_sample_req
      -- CP-element group 199: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_loopback_sample_req_ps
      -- 
    phi_stmt_589_loopback_sample_req_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_loopback_sample_req_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(199), ack => phi_stmt_589_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(199) is bound as output of CP function.
    -- CP-element group 200:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	130 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_entry_trigger
      -- 
    zeropad_same_CP_159_elements(200) <= zeropad_same_CP_159_elements(130);
    -- CP-element group 201:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_entry_sample_req
      -- CP-element group 201: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_entry_sample_req_ps
      -- 
    phi_stmt_589_entry_sample_req_1349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_entry_sample_req_1349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(201), ack => phi_stmt_589_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(201) is bound as output of CP function.
    -- CP-element group 202:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_phi_mux_ack_ps
      -- CP-element group 202: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_589_phi_mux_ack
      -- 
    phi_stmt_589_phi_mux_ack_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_589_ack_0, ack => zeropad_same_CP_159_elements(202)); -- 
    -- CP-element group 203:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (4) 
      -- CP-element group 203: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_sample_start__ps
      -- CP-element group 203: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Sample/req
      -- 
    req_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(203), ack => add_dest_dim0_init_567_591_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(203) is bound as output of CP function.
    -- CP-element group 204:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (4) 
      -- CP-element group 204: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_update_start__ps
      -- CP-element group 204: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_update_start_
      -- CP-element group 204: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Update/req
      -- 
    req_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(204), ack => add_dest_dim0_init_567_591_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(204) is bound as output of CP function.
    -- CP-element group 205:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (4) 
      -- CP-element group 205: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_sample_completed__ps
      -- CP-element group 205: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Sample/ack
      -- 
    ack_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_567_591_buf_ack_0, ack => zeropad_same_CP_159_elements(205)); -- 
    -- CP-element group 206:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (4) 
      -- CP-element group 206: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_update_completed__ps
      -- CP-element group 206: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim0_init_591_Update/ack
      -- 
    ack_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_567_591_buf_ack_1, ack => zeropad_same_CP_159_elements(206)); -- 
    -- CP-element group 207:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (4) 
      -- CP-element group 207: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_sample_start__ps
      -- CP-element group 207: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Sample/req
      -- 
    req_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(207), ack => next_add_dest_dim0_734_592_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(207) is bound as output of CP function.
    -- CP-element group 208:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (4) 
      -- CP-element group 208: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_update_start__ps
      -- CP-element group 208: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_update_start_
      -- CP-element group 208: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Update/req
      -- 
    req_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(208), ack => next_add_dest_dim0_734_592_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(208) is bound as output of CP function.
    -- CP-element group 209:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (4) 
      -- CP-element group 209: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_sample_completed__ps
      -- CP-element group 209: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Sample/ack
      -- 
    ack_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_734_592_buf_ack_0, ack => zeropad_same_CP_159_elements(209)); -- 
    -- CP-element group 210:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (4) 
      -- CP-element group 210: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_update_completed__ps
      -- CP-element group 210: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim0_592_Update/ack
      -- 
    ack_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_734_592_buf_ack_1, ack => zeropad_same_CP_159_elements(210)); -- 
    -- CP-element group 211:  join  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	131 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	134 
    -- CP-element group 211: 	279 
    -- CP-element group 211: 	283 
    -- CP-element group 211: 	287 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	133 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_sample_start_
      -- 
    zeropad_same_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(279) & zeropad_same_CP_159_elements(283) & zeropad_same_CP_159_elements(287);
      gj_zeropad_same_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	131 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	216 
    -- CP-element group 212: 	264 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	135 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_update_start_
      -- 
    zeropad_same_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(216) & zeropad_same_CP_159_elements(264);
      gj_zeropad_same_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	133 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_sample_start__ps
      -- 
    zeropad_same_CP_159_elements(213) <= zeropad_same_CP_159_elements(133);
    -- CP-element group 214:  join  transition  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	134 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(214) is bound as output of CP function.
    -- CP-element group 215:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	135 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_update_start__ps
      -- 
    zeropad_same_CP_159_elements(215) <= zeropad_same_CP_159_elements(135);
    -- CP-element group 216:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	136 
    -- CP-element group 216: 	262 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	212 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_update_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(216) is bound as output of CP function.
    -- CP-element group 217:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	129 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_loopback_trigger
      -- 
    zeropad_same_CP_159_elements(217) <= zeropad_same_CP_159_elements(129);
    -- CP-element group 218:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_loopback_sample_req
      -- CP-element group 218: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_loopback_sample_req_ps
      -- 
    phi_stmt_593_loopback_sample_req_1400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_593_loopback_sample_req_1400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(218), ack => phi_stmt_593_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(218) is bound as output of CP function.
    -- CP-element group 219:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	130 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_entry_trigger
      -- 
    zeropad_same_CP_159_elements(219) <= zeropad_same_CP_159_elements(130);
    -- CP-element group 220:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_entry_sample_req
      -- CP-element group 220: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_entry_sample_req_ps
      -- 
    phi_stmt_593_entry_sample_req_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_593_entry_sample_req_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(220), ack => phi_stmt_593_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(220) is bound as output of CP function.
    -- CP-element group 221:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_phi_mux_ack
      -- CP-element group 221: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_593_phi_mux_ack_ps
      -- 
    phi_stmt_593_phi_mux_ack_1406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_593_ack_0, ack => zeropad_same_CP_159_elements(221)); -- 
    -- CP-element group 222:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (4) 
      -- CP-element group 222: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_sample_start__ps
      -- CP-element group 222: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Sample/req
      -- 
    req_1419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(222), ack => add_dest_dim1_init_570_595_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(222) is bound as output of CP function.
    -- CP-element group 223:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (4) 
      -- CP-element group 223: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_update_start__ps
      -- CP-element group 223: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_update_start_
      -- CP-element group 223: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Update/req
      -- 
    req_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(223), ack => add_dest_dim1_init_570_595_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(223) is bound as output of CP function.
    -- CP-element group 224:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (4) 
      -- CP-element group 224: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_sample_completed__ps
      -- CP-element group 224: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Sample/ack
      -- 
    ack_1420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_570_595_buf_ack_0, ack => zeropad_same_CP_159_elements(224)); -- 
    -- CP-element group 225:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (4) 
      -- CP-element group 225: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_update_completed__ps
      -- CP-element group 225: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_dest_dim1_init_595_Update/ack
      -- 
    ack_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_570_595_buf_ack_1, ack => zeropad_same_CP_159_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_sample_start__ps
      -- CP-element group 226: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Sample/req
      -- 
    req_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(226), ack => next_add_dest_dim1_728_596_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(226) is bound as output of CP function.
    -- CP-element group 227:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_update_start__ps
      -- CP-element group 227: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_update_start_
      -- CP-element group 227: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Update/req
      -- 
    req_1442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(227), ack => next_add_dest_dim1_728_596_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(227) is bound as output of CP function.
    -- CP-element group 228:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (4) 
      -- CP-element group 228: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_sample_completed__ps
      -- CP-element group 228: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Sample/ack
      -- 
    ack_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_728_596_buf_ack_0, ack => zeropad_same_CP_159_elements(228)); -- 
    -- CP-element group 229:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (4) 
      -- CP-element group 229: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_update_completed__ps
      -- CP-element group 229: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_dest_dim1_596_Update/ack
      -- 
    ack_1443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_728_596_buf_ack_1, ack => zeropad_same_CP_159_elements(229)); -- 
    -- CP-element group 230:  join  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	131 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	134 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	133 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_sample_start_
      -- 
    zeropad_same_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(134);
      gj_zeropad_same_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	131 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	235 
    -- CP-element group 231: 	252 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	135 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_update_start_
      -- 
    zeropad_same_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(235) & zeropad_same_CP_159_elements(252);
      gj_zeropad_same_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	133 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_sample_start__ps
      -- 
    zeropad_same_CP_159_elements(232) <= zeropad_same_CP_159_elements(133);
    -- CP-element group 233:  join  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	134 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_159_elements(233) is bound as output of CP function.
    -- CP-element group 234:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	135 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_update_start__ps
      -- 
    zeropad_same_CP_159_elements(234) <= zeropad_same_CP_159_elements(135);
    -- CP-element group 235:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	136 
    -- CP-element group 235: 	252 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	231 
    -- CP-element group 235:  members (15) 
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_update_completed__ps
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_resized_1
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_scaled_1
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_computed_1
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_resize_1/$entry
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_resize_1/$exit
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_resize_1/index_resize_req
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_resize_1/index_resize_ack
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_scale_1/$entry
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_scale_1/$exit
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_scale_1/scale_rename_req
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_index_scale_1/scale_rename_ack
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Sample/req
      -- 
    req_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(235), ack => array_obj_ref_632_index_offset_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(235) is bound as output of CP function.
    -- CP-element group 236:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	129 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_loopback_trigger
      -- 
    zeropad_same_CP_159_elements(236) <= zeropad_same_CP_159_elements(129);
    -- CP-element group 237:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_loopback_sample_req
      -- CP-element group 237: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_loopback_sample_req_ps
      -- 
    phi_stmt_597_loopback_sample_req_1454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_597_loopback_sample_req_1454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(237), ack => phi_stmt_597_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(237) is bound as output of CP function.
    -- CP-element group 238:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	130 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_entry_trigger
      -- 
    zeropad_same_CP_159_elements(238) <= zeropad_same_CP_159_elements(130);
    -- CP-element group 239:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_entry_sample_req
      -- CP-element group 239: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_entry_sample_req_ps
      -- 
    phi_stmt_597_entry_sample_req_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_597_entry_sample_req_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(239), ack => phi_stmt_597_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(239) is bound as output of CP function.
    -- CP-element group 240:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_phi_mux_ack
      -- CP-element group 240: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/phi_stmt_597_phi_mux_ack_ps
      -- 
    phi_stmt_597_phi_mux_ack_1460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_597_ack_0, ack => zeropad_same_CP_159_elements(240)); -- 
    -- CP-element group 241:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_sample_start__ps
      -- CP-element group 241: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_sample_completed__ps
      -- CP-element group 241: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_sample_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(241) is bound as output of CP function.
    -- CP-element group 242:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_update_start__ps
      -- CP-element group 242: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_update_start_
      -- 
    -- Element group zeropad_same_CP_159_elements(242) is bound as output of CP function.
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_update_completed__ps
      -- 
    zeropad_same_CP_159_elements(243) <= zeropad_same_CP_159_elements(244);
    -- CP-element group 244:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	243 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_add_src_init_599_update_completed_
      -- 
    -- Element group zeropad_same_CP_159_elements(244) is a control-delay.
    cp_element_244_delay: control_delay_element  generic map(name => " 244_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(242), ack => zeropad_same_CP_159_elements(244), clk => clk, reset =>reset);
    -- CP-element group 245:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_sample_start__ps
      -- CP-element group 245: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Sample/req
      -- 
    req_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(245), ack => next_add_src_715_600_buf_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(245) is bound as output of CP function.
    -- CP-element group 246:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_update_start__ps
      -- CP-element group 246: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_update_start_
      -- CP-element group 246: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Update/req
      -- 
    req_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(246), ack => next_add_src_715_600_buf_req_1); -- 
    -- Element group zeropad_same_CP_159_elements(246) is bound as output of CP function.
    -- CP-element group 247:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (4) 
      -- CP-element group 247: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_sample_completed__ps
      -- CP-element group 247: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Sample/ack
      -- 
    ack_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_715_600_buf_ack_0, ack => zeropad_same_CP_159_elements(247)); -- 
    -- CP-element group 248:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (4) 
      -- CP-element group 248: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_update_completed__ps
      -- CP-element group 248: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/R_next_add_src_600_Update/ack
      -- 
    ack_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_715_600_buf_ack_1, ack => zeropad_same_CP_159_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	253 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	254 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	254 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_request/$entry
      -- CP-element group 249: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_request/req
      -- 
    req_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(249), ack => addr_of_633_final_reg_req_0); -- 
    zeropad_same_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(253) & zeropad_same_CP_159_elements(254);
      gj_zeropad_same_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	131 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	255 
    -- CP-element group 250: 	258 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	255 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_update_start_
      -- CP-element group 250: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_complete/$entry
      -- CP-element group 250: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_complete/req
      -- 
    req_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(250), ack => addr_of_633_final_reg_req_1); -- 
    zeropad_same_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(255) & zeropad_same_CP_159_elements(258);
      gj_zeropad_same_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	131 
    -- CP-element group 251: marked-predecessors 
    -- CP-element group 251: 	253 
    -- CP-element group 251: 	254 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_update_start
      -- CP-element group 251: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Update/req
      -- 
    req_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(251), ack => array_obj_ref_632_index_offset_req_1); -- 
    zeropad_same_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(253) & zeropad_same_CP_159_elements(254);
      gj_zeropad_same_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	235 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	293 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	231 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_sample_complete
      -- CP-element group 252: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Sample/ack
      -- 
    ack_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_632_index_offset_ack_0, ack => zeropad_same_CP_159_elements(252)); -- 
    -- CP-element group 253:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	249 
    -- CP-element group 253: marked-successors 
    -- CP-element group 253: 	251 
    -- CP-element group 253:  members (8) 
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_root_address_calculated
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_offset_calculated
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_final_index_sum_regn_Update/ack
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_base_plus_offset/$entry
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_base_plus_offset/$exit
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_base_plus_offset/sum_rename_req
      -- CP-element group 253: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_632_base_plus_offset/sum_rename_ack
      -- 
    ack_1519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_632_index_offset_ack_1, ack => zeropad_same_CP_159_elements(253)); -- 
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	249 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	249 
    -- CP-element group 254: 	251 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_request/$exit
      -- CP-element group 254: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_request/ack
      -- 
    ack_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_633_final_reg_ack_0, ack => zeropad_same_CP_159_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	250 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	250 
    -- CP-element group 255:  members (19) 
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_complete/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_633_complete/ack
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_address_calculated
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_word_address_calculated
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_root_address_calculated
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_address_resized
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_addr_resize/$entry
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_addr_resize/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_addr_resize/base_resize_req
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_addr_resize/base_resize_ack
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_plus_offset/$entry
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_plus_offset/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_plus_offset/sum_rename_req
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_base_plus_offset/sum_rename_ack
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_word_addrgen/$entry
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_word_addrgen/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_word_addrgen/root_register_req
      -- CP-element group 255: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_word_addrgen/root_register_ack
      -- 
    ack_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_633_final_reg_ack_1, ack => zeropad_same_CP_159_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (5) 
      -- CP-element group 256: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/word_access_start/$entry
      -- CP-element group 256: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/word_access_start/word_0/$entry
      -- CP-element group 256: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/word_access_start/word_0/rr
      -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(256), ack => ptr_deref_637_load_0_req_0); -- 
    zeropad_same_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(255) & zeropad_same_CP_159_elements(258);
      gj_zeropad_same_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: 	274 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (5) 
      -- CP-element group 257: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_update_start_
      -- CP-element group 257: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/word_access_complete/$entry
      -- CP-element group 257: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/word_access_complete/word_0/$entry
      -- CP-element group 257: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/word_access_complete/word_0/cr
      -- 
    cr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(257), ack => ptr_deref_637_load_0_req_1); -- 
    zeropad_same_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(259) & zeropad_same_CP_159_elements(274);
      gj_zeropad_same_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	250 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (5) 
      -- CP-element group 258: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/word_access_start/$exit
      -- CP-element group 258: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/word_access_start/word_0/$exit
      -- CP-element group 258: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Sample/word_access_start/word_0/ra
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_637_load_0_ack_0, ack => zeropad_same_CP_159_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	272 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (9) 
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/word_access_complete/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/word_access_complete/word_0/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/word_access_complete/word_0/ca
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/ptr_deref_637_Merge/$entry
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/ptr_deref_637_Merge/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/ptr_deref_637_Merge/merge_req
      -- CP-element group 259: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_637_Update/ptr_deref_637_Merge/merge_ack
      -- 
    ca_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_637_load_0_ack_1, ack => zeropad_same_CP_159_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	265 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	266 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	266 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_request/$entry
      -- CP-element group 260: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_request/req
      -- 
    req_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(260), ack => addr_of_645_final_reg_req_0); -- 
    zeropad_same_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(265) & zeropad_same_CP_159_elements(266);
      gj_zeropad_same_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	131 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	267 
    -- CP-element group 261: 	270 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	267 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_update_start_
      -- CP-element group 261: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_complete/$entry
      -- CP-element group 261: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_complete/req
      -- 
    req_1629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(261), ack => addr_of_645_final_reg_req_1); -- 
    zeropad_same_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(267) & zeropad_same_CP_159_elements(270);
      gj_zeropad_same_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	178 
    -- CP-element group 262: 	197 
    -- CP-element group 262: 	216 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (13) 
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_resized_1
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_scaled_1
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_computed_1
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_resize_1/$entry
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_resize_1/$exit
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_resize_1/index_resize_req
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_resize_1/index_resize_ack
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_scale_1/$entry
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_scale_1/$exit
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_scale_1/scale_rename_req
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_index_scale_1/scale_rename_ack
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Sample/req
      -- 
    req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(262), ack => array_obj_ref_644_index_offset_req_0); -- 
    zeropad_same_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(178) & zeropad_same_CP_159_elements(197) & zeropad_same_CP_159_elements(216);
      gj_zeropad_same_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	131 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: 	266 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_update_start
      -- CP-element group 263: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Update/req
      -- 
    req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(263), ack => array_obj_ref_644_index_offset_req_1); -- 
    zeropad_same_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(265) & zeropad_same_CP_159_elements(266);
      gj_zeropad_same_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	293 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	174 
    -- CP-element group 264: 	193 
    -- CP-element group 264: 	212 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_sample_complete
      -- CP-element group 264: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Sample/ack
      -- 
    ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_644_index_offset_ack_0, ack => zeropad_same_CP_159_elements(264)); -- 
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	260 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (8) 
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_root_address_calculated
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_offset_calculated
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_final_index_sum_regn_Update/ack
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_base_plus_offset/$entry
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_base_plus_offset/$exit
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_base_plus_offset/sum_rename_req
      -- CP-element group 265: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/array_obj_ref_644_base_plus_offset/sum_rename_ack
      -- 
    ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_644_index_offset_ack_1, ack => zeropad_same_CP_159_elements(265)); -- 
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	260 
    -- CP-element group 266: successors 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	260 
    -- CP-element group 266: 	263 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_request/$exit
      -- CP-element group 266: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_request/ack
      -- 
    ack_1625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_645_final_reg_ack_0, ack => zeropad_same_CP_159_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	261 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	261 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_complete/$exit
      -- CP-element group 267: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/addr_of_645_complete/ack
      -- 
    ack_1630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_645_final_reg_ack_1, ack => zeropad_same_CP_159_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Sample/req
      -- 
    req_1638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(268), ack => W_ov_647_delayed_6_0_647_inst_req_0); -- 
    zeropad_same_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(267) & zeropad_same_CP_159_elements(270);
      gj_zeropad_same_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	274 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_update_start_
      -- CP-element group 269: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Update/req
      -- 
    req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(269), ack => W_ov_647_delayed_6_0_647_inst_req_1); -- 
    zeropad_same_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(271) & zeropad_same_CP_159_elements(274);
      gj_zeropad_same_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	261 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Sample/ack
      -- 
    ack_1639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ov_647_delayed_6_0_647_inst_ack_0, ack => zeropad_same_CP_159_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (19) 
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_649_Update/ack
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_address_calculated
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_word_address_calculated
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_root_address_calculated
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_address_resized
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_addr_resize/$entry
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_addr_resize/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_addr_resize/base_resize_req
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_addr_resize/base_resize_ack
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_plus_offset/$entry
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_plus_offset/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_plus_offset/sum_rename_req
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_base_plus_offset/sum_rename_ack
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_word_addrgen/$entry
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_word_addrgen/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_word_addrgen/root_register_req
      -- CP-element group 271: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_word_addrgen/root_register_ack
      -- 
    ack_1644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ov_647_delayed_6_0_647_inst_ack_1, ack => zeropad_same_CP_159_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	259 
    -- CP-element group 272: 	271 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (9) 
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/ptr_deref_651_Split/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/ptr_deref_651_Split/$exit
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/ptr_deref_651_Split/split_req
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/ptr_deref_651_Split/split_ack
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/word_access_start/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/word_access_start/word_0/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/word_access_start/word_0/rr
      -- 
    rr_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(272), ack => ptr_deref_651_store_0_req_0); -- 
    zeropad_same_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(259) & zeropad_same_CP_159_elements(271) & zeropad_same_CP_159_elements(274);
      gj_zeropad_same_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (5) 
      -- CP-element group 273: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_update_start_
      -- CP-element group 273: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/word_access_complete/$entry
      -- CP-element group 273: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/word_access_complete/word_0/$entry
      -- CP-element group 273: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/word_access_complete/word_0/cr
      -- 
    cr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(273), ack => ptr_deref_651_store_0_req_1); -- 
    zeropad_same_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_same_CP_159_elements(275);
      gj_zeropad_same_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	257 
    -- CP-element group 274: 	269 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (5) 
      -- CP-element group 274: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/word_access_start/$exit
      -- CP-element group 274: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/word_access_start/word_0/$exit
      -- CP-element group 274: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Sample/word_access_start/word_0/ra
      -- 
    ra_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_651_store_0_ack_0, ack => zeropad_same_CP_159_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	293 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (5) 
      -- CP-element group 275: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/word_access_complete/$exit
      -- CP-element group 275: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/word_access_complete/word_0/$exit
      -- CP-element group 275: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/ptr_deref_651_Update/word_access_complete/word_0/ca
      -- 
    ca_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_651_store_0_ack_1, ack => zeropad_same_CP_159_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	131 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Sample/req
      -- 
    req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(276), ack => W_dim2_limit_658_delayed_1_0_659_inst_req_0); -- 
    zeropad_same_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(278);
      gj_zeropad_same_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	134 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_update_start_
      -- CP-element group 277: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Update/req
      -- 
    req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(277), ack => W_dim2_limit_658_delayed_1_0_659_inst_req_1); -- 
    zeropad_same_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(279);
      gj_zeropad_same_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Sample/ack
      -- 
    ack_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_658_delayed_1_0_659_inst_ack_0, ack => zeropad_same_CP_159_elements(278)); -- 
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	132 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	137 
    -- CP-element group 279: 	154 
    -- CP-element group 279: 	173 
    -- CP-element group 279: 	192 
    -- CP-element group 279: 	211 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_661_Update/ack
      -- 
    ack_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_658_delayed_1_0_659_inst_ack_1, ack => zeropad_same_CP_159_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	131 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Sample/rr
      -- 
    rr_1716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(280), ack => SUB_u16_u16_670_inst_req_0); -- 
    zeropad_same_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(282);
      gj_zeropad_same_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	134 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_update_start_
      -- CP-element group 281: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Update/cr
      -- 
    cr_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(281), ack => SUB_u16_u16_670_inst_req_1); -- 
    zeropad_same_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(283);
      gj_zeropad_same_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Sample/ra
      -- 
    ra_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_670_inst_ack_0, ack => zeropad_same_CP_159_elements(282)); -- 
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	132 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	137 
    -- CP-element group 283: 	154 
    -- CP-element group 283: 	192 
    -- CP-element group 283: 	211 
    -- CP-element group 283: 	281 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_670_Update/ca
      -- 
    ca_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_670_inst_ack_1, ack => zeropad_same_CP_159_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	131 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Sample/req
      -- 
    req_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(284), ack => W_nid1_true4_711_delayed_1_0_716_inst_req_0); -- 
    zeropad_same_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(286);
      gj_zeropad_same_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	134 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_update_start_
      -- CP-element group 285: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Update/req
      -- 
    req_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(285), ack => W_nid1_true4_711_delayed_1_0_716_inst_req_1); -- 
    zeropad_same_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(287);
      gj_zeropad_same_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Sample/ack
      -- 
    ack_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true4_711_delayed_1_0_716_inst_ack_0, ack => zeropad_same_CP_159_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	293 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	211 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/assign_stmt_718_Update/ack
      -- 
    ack_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true4_711_delayed_1_0_716_inst_ack_1, ack => zeropad_same_CP_159_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	131 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Sample/rr
      -- 
    rr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(288), ack => SUB_u16_u16_760_inst_req_0); -- 
    zeropad_same_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(131) & zeropad_same_CP_159_elements(290);
      gj_zeropad_same_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_update_start_
      -- CP-element group 289: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Update/cr
      -- 
    cr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(289), ack => SUB_u16_u16_760_inst_req_1); -- 
    zeropad_same_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_same_CP_159_elements(291);
      gj_zeropad_same_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Sample/ra
      -- 
    ra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_760_inst_ack_0, ack => zeropad_same_CP_159_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	132 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/SUB_u16_u16_760_Update/ca
      -- 
    ca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_760_inst_ack_1, ack => zeropad_same_CP_159_elements(291)); -- 
    -- CP-element group 292:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	131 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	132 
    -- CP-element group 292:  members (1) 
      -- CP-element group 292: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group zeropad_same_CP_159_elements(292) is a control-delay.
    cp_element_292_delay: control_delay_element  generic map(name => " 292_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(131), ack => zeropad_same_CP_159_elements(292), clk => clk, reset =>reset);
    -- CP-element group 293:  join  transition  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	134 
    -- CP-element group 293: 	252 
    -- CP-element group 293: 	264 
    -- CP-element group 293: 	275 
    -- CP-element group 293: 	287 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	128 
    -- CP-element group 293:  members (1) 
      -- CP-element group 293: 	 branch_block_stmt_38/do_while_stmt_575/do_while_stmt_575_loop_body/$exit
      -- 
    zeropad_same_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(134) & zeropad_same_CP_159_elements(252) & zeropad_same_CP_159_elements(264) & zeropad_same_CP_159_elements(275) & zeropad_same_CP_159_elements(287);
      gj_zeropad_same_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	127 
    -- CP-element group 294: successors 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_38/do_while_stmt_575/loop_exit/$exit
      -- CP-element group 294: 	 branch_block_stmt_38/do_while_stmt_575/loop_exit/ack
      -- 
    ack_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_575_branch_ack_0, ack => zeropad_same_CP_159_elements(294)); -- 
    -- CP-element group 295:  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	127 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (2) 
      -- CP-element group 295: 	 branch_block_stmt_38/do_while_stmt_575/loop_taken/$exit
      -- CP-element group 295: 	 branch_block_stmt_38/do_while_stmt_575/loop_taken/ack
      -- 
    ack_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_575_branch_ack_1, ack => zeropad_same_CP_159_elements(295)); -- 
    -- CP-element group 296:  transition  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	125 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	1 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_38/do_while_stmt_575/$exit
      -- 
    zeropad_same_CP_159_elements(296) <= zeropad_same_CP_159_elements(125);
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	1 
    -- CP-element group 297: successors 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Sample/cra
      -- CP-element group 297: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Sample/$exit
      -- 
    cra_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_777_call_ack_0, ack => zeropad_same_CP_159_elements(297)); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	1 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	301 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_Update/cca
      -- CP-element group 298: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/call_stmt_777_update_completed_
      -- 
    cca_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_777_call_ack_1, ack => zeropad_same_CP_159_elements(298)); -- 
    rr_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(298), ack => type_cast_787_inst_req_0); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	1 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Sample/ra
      -- CP-element group 299: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Sample/$exit
      -- 
    ra_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_0, ack => zeropad_same_CP_159_elements(299)); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	1 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	303 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_782_Update/ca
      -- 
    ca_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_1, ack => zeropad_same_CP_159_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	298 
    -- CP-element group 301: successors 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Sample/ra
      -- CP-element group 301: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Sample/$exit
      -- 
    ra_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_0, ack => zeropad_same_CP_159_elements(301)); -- 
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	1 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Update/ca
      -- CP-element group 302: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/type_cast_787_update_completed_
      -- 
    ca_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_1, ack => zeropad_same_CP_159_elements(302)); -- 
    -- CP-element group 303:  join  fork  transition  place  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	300 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303: 	305 
    -- CP-element group 303: 	306 
    -- CP-element group 303: 	307 
    -- CP-element group 303: 	308 
    -- CP-element group 303: 	309 
    -- CP-element group 303: 	310 
    -- CP-element group 303: 	311 
    -- CP-element group 303: 	312 
    -- CP-element group 303: 	313 
    -- CP-element group 303: 	314 
    -- CP-element group 303: 	315 
    -- CP-element group 303: 	316 
    -- CP-element group 303: 	317 
    -- CP-element group 303: 	318 
    -- CP-element group 303: 	319 
    -- CP-element group 303:  members (52) 
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793__exit__
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892__entry__
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Update/cr
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/call_stmt_777_to_assign_stmt_793/$exit
      -- 
    rr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_837_inst_req_0); -- 
    rr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_797_inst_req_0); -- 
    rr_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_817_inst_req_0); -- 
    cr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_837_inst_req_1); -- 
    cr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_797_inst_req_1); -- 
    cr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_817_inst_req_1); -- 
    rr_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_827_inst_req_0); -- 
    rr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_847_inst_req_0); -- 
    cr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_827_inst_req_1); -- 
    cr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_807_inst_req_1); -- 
    cr_1919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_867_inst_req_1); -- 
    rr_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_867_inst_req_0); -- 
    rr_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_807_inst_req_0); -- 
    cr_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_857_inst_req_1); -- 
    rr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_857_inst_req_0); -- 
    cr_1891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(303), ack => type_cast_847_inst_req_1); -- 
    zeropad_same_cp_element_group_303: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_303"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(300) & zeropad_same_CP_159_elements(302);
      gj_zeropad_same_cp_element_group_303 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(303), clk => clk, reset => reset); --
    end block;
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_sample_completed_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Sample/ra
      -- 
    ra_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_0, ack => zeropad_same_CP_159_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	303 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	340 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_update_completed_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_797_Update/ca
      -- 
    ca_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_1, ack => zeropad_same_CP_159_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	303 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Sample/ra
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_sample_completed_
      -- 
    ra_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_0, ack => zeropad_same_CP_159_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	303 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	337 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Update/ca
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_807_update_completed_
      -- 
    ca_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_1, ack => zeropad_same_CP_159_elements(307)); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	303 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Sample/$exit
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Sample/ra
      -- 
    ra_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => zeropad_same_CP_159_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	303 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	334 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_update_completed_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_817_Update/ca
      -- 
    ca_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => zeropad_same_CP_159_elements(309)); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	303 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Sample/ra
      -- 
    ra_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_0, ack => zeropad_same_CP_159_elements(310)); -- 
    -- CP-element group 311:  transition  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	303 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	331 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_827_Update/ca
      -- 
    ca_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_1, ack => zeropad_same_CP_159_elements(311)); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	303 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Sample/ra
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Sample/$exit
      -- 
    ra_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_0, ack => zeropad_same_CP_159_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	303 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	328 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_837_Update/ca
      -- 
    ca_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_1, ack => zeropad_same_CP_159_elements(313)); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	303 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Sample/ra
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Sample/$exit
      -- 
    ra_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => zeropad_same_CP_159_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	303 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	325 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Update/ca
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_847_Update/$exit
      -- 
    ca_1892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_1, ack => zeropad_same_CP_159_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	303 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Sample/ra
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_sample_completed_
      -- 
    ra_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_0, ack => zeropad_same_CP_159_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	303 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	322 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Update/ca
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_857_update_completed_
      -- 
    ca_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_1, ack => zeropad_same_CP_159_elements(317)); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	303 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Sample/ra
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_sample_completed_
      -- 
    ra_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_867_inst_ack_0, ack => zeropad_same_CP_159_elements(318)); -- 
    -- CP-element group 319:  transition  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	303 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (6) 
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Sample/req
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_sample_start_
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Update/ca
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/type_cast_867_update_completed_
      -- 
    ca_1920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_867_inst_ack_1, ack => zeropad_same_CP_159_elements(319)); -- 
    req_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(319), ack => WPIPE_ConvTranspose_output_pipe_869_inst_req_0); -- 
    -- CP-element group 320:  transition  input  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (6) 
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Update/req
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Update/$entry
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Sample/ack
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_update_start_
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_sample_completed_
      -- 
    ack_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_869_inst_ack_0, ack => zeropad_same_CP_159_elements(320)); -- 
    req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(320), ack => WPIPE_ConvTranspose_output_pipe_869_inst_req_1); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Update/ack
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_869_update_completed_
      -- 
    ack_1934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_869_inst_ack_1, ack => zeropad_same_CP_159_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	317 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Sample/req
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_sample_start_
      -- 
    req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(322), ack => WPIPE_ConvTranspose_output_pipe_872_inst_req_0); -- 
    zeropad_same_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(317) & zeropad_same_CP_159_elements(321);
      gj_zeropad_same_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Update/req
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_update_start_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_sample_completed_
      -- 
    ack_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_872_inst_ack_0, ack => zeropad_same_CP_159_elements(323)); -- 
    req_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(323), ack => WPIPE_ConvTranspose_output_pipe_872_inst_req_1); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_872_update_completed_
      -- 
    ack_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_872_inst_ack_1, ack => zeropad_same_CP_159_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	315 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Sample/req
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_sample_start_
      -- 
    req_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(325), ack => WPIPE_ConvTranspose_output_pipe_875_inst_req_0); -- 
    zeropad_same_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(315) & zeropad_same_CP_159_elements(324);
      gj_zeropad_same_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Update/req
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Sample/ack
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Sample/$exit
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_update_start_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_sample_completed_
      -- 
    ack_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_875_inst_ack_0, ack => zeropad_same_CP_159_elements(326)); -- 
    req_1961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(326), ack => WPIPE_ConvTranspose_output_pipe_875_inst_req_1); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Update/ack
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_Update/$exit
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_875_update_completed_
      -- 
    ack_1962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_875_inst_ack_1, ack => zeropad_same_CP_159_elements(327)); -- 
    -- CP-element group 328:  join  transition  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	313 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Sample/req
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_sample_start_
      -- 
    req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(328), ack => WPIPE_ConvTranspose_output_pipe_878_inst_req_0); -- 
    zeropad_same_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(313) & zeropad_same_CP_159_elements(327);
      gj_zeropad_same_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Update/req
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_update_start_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_sample_completed_
      -- 
    ack_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_878_inst_ack_0, ack => zeropad_same_CP_159_elements(329)); -- 
    req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(329), ack => WPIPE_ConvTranspose_output_pipe_878_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_878_Update/ack
      -- 
    ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_878_inst_ack_1, ack => zeropad_same_CP_159_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	311 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Sample/req
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_sample_start_
      -- 
    req_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(331), ack => WPIPE_ConvTranspose_output_pipe_881_inst_req_0); -- 
    zeropad_same_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(311) & zeropad_same_CP_159_elements(330);
      gj_zeropad_same_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_update_start_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Sample/ack
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Update/$entry
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Update/req
      -- 
    ack_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_881_inst_ack_0, ack => zeropad_same_CP_159_elements(332)); -- 
    req_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(332), ack => WPIPE_ConvTranspose_output_pipe_881_inst_req_1); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_881_Update/ack
      -- 
    ack_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_881_inst_ack_1, ack => zeropad_same_CP_159_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	309 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Sample/req
      -- 
    req_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(334), ack => WPIPE_ConvTranspose_output_pipe_884_inst_req_0); -- 
    zeropad_same_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(309) & zeropad_same_CP_159_elements(333);
      gj_zeropad_same_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_update_start_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Update/req
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Update/$entry
      -- 
    ack_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_884_inst_ack_0, ack => zeropad_same_CP_159_elements(335)); -- 
    req_2003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(335), ack => WPIPE_ConvTranspose_output_pipe_884_inst_req_1); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_884_Update/$exit
      -- 
    ack_2004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_884_inst_ack_1, ack => zeropad_same_CP_159_elements(336)); -- 
    -- CP-element group 337:  join  transition  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	307 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Sample/req
      -- 
    req_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(337), ack => WPIPE_ConvTranspose_output_pipe_887_inst_req_0); -- 
    zeropad_same_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(307) & zeropad_same_CP_159_elements(336);
      gj_zeropad_same_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Update/req
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_sample_completed_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_update_start_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Sample/ack
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Update/$entry
      -- 
    ack_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_887_inst_ack_0, ack => zeropad_same_CP_159_elements(338)); -- 
    req_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(338), ack => WPIPE_ConvTranspose_output_pipe_887_inst_req_1); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Update/ack
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_update_completed_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_887_Update/$exit
      -- 
    ack_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_887_inst_ack_1, ack => zeropad_same_CP_159_elements(339)); -- 
    -- CP-element group 340:  join  transition  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	305 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Sample/req
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_sample_start_
      -- 
    req_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(340), ack => WPIPE_ConvTranspose_output_pipe_890_inst_req_0); -- 
    zeropad_same_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(305) & zeropad_same_CP_159_elements(339);
      gj_zeropad_same_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Update/req
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_update_start_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_sample_completed_
      -- 
    ack_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_890_inst_ack_0, ack => zeropad_same_CP_159_elements(341)); -- 
    req_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(341), ack => WPIPE_ConvTranspose_output_pipe_890_inst_req_1); -- 
    -- CP-element group 342:  branch  transition  place  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (17) 
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900_if_link/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_899/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/R_cmp264449_901_place
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900_dead_link/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892__exit__
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_899__entry__
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_899__exit__
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900__entry__
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_798_to_assign_stmt_892/WPIPE_ConvTranspose_output_pipe_890_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_899/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900_eval_test/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900_eval_test/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900_eval_test/branch_req
      -- CP-element group 342: 	 branch_block_stmt_38/if_stmt_900_else_link/$entry
      -- 
    ack_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_890_inst_ack_1, ack => zeropad_same_CP_159_elements(342)); -- 
    branch_req_2043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(342), ack => if_stmt_900_branch_req_0); -- 
    -- CP-element group 343:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343: 	346 
    -- CP-element group 343:  members (18) 
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_sample_start_
      -- CP-element group 343: 	 branch_block_stmt_38/merge_stmt_906__exit__
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941__entry__
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_update_start_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Sample/rr
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/forx_xend273_bbx_xnph
      -- CP-element group 343: 	 branch_block_stmt_38/if_stmt_900_if_link/if_choice_transition
      -- CP-element group 343: 	 branch_block_stmt_38/if_stmt_900_if_link/$exit
      -- CP-element group 343: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 343: 	 branch_block_stmt_38/merge_stmt_906_PhiReqMerge
      -- CP-element group 343: 	 branch_block_stmt_38/merge_stmt_906_PhiAck/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/merge_stmt_906_PhiAck/$exit
      -- CP-element group 343: 	 branch_block_stmt_38/merge_stmt_906_PhiAck/dummy
      -- 
    if_choice_transition_2048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_900_branch_ack_1, ack => zeropad_same_CP_159_elements(343)); -- 
    rr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(343), ack => type_cast_927_inst_req_0); -- 
    cr_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(343), ack => type_cast_927_inst_req_1); -- 
    -- CP-element group 344:  transition  place  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	415 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 branch_block_stmt_38/forx_xend273_forx_xend444
      -- CP-element group 344: 	 branch_block_stmt_38/if_stmt_900_else_link/else_choice_transition
      -- CP-element group 344: 	 branch_block_stmt_38/if_stmt_900_else_link/$exit
      -- CP-element group 344: 	 branch_block_stmt_38/forx_xend273_forx_xend444_PhiReq/$entry
      -- CP-element group 344: 	 branch_block_stmt_38/forx_xend273_forx_xend444_PhiReq/$exit
      -- 
    else_choice_transition_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_900_branch_ack_0, ack => zeropad_same_CP_159_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Sample/ra
      -- 
    ra_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => zeropad_same_CP_159_elements(345)); -- 
    -- CP-element group 346:  transition  place  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	343 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	409 
    -- CP-element group 346:  members (9) 
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/$exit
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941__exit__
      -- CP-element group 346: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_912_to_assign_stmt_941/type_cast_927_Update/ca
      -- CP-element group 346: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_944/$entry
      -- CP-element group 346: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/$entry
      -- 
    ca_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => zeropad_same_CP_159_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	414 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	392 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_sample_complete
      -- 
    ack_2100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_offset_ack_0, ack => zeropad_same_CP_159_elements(347)); -- 
    -- CP-element group 348:  transition  input  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	414 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (11) 
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_root_address_calculated
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_offset_calculated
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_request/req
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_request/$entry
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_base_plus_offset/sum_rename_ack
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_base_plus_offset/sum_rename_req
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Update/ack
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_base_plus_offset/$entry
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_base_plus_offset/$exit
      -- 
    ack_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_offset_ack_1, ack => zeropad_same_CP_159_elements(348)); -- 
    req_2114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(348), ack => addr_of_957_final_reg_req_0); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_request/ack
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_request/$exit
      -- 
    ack_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_957_final_reg_ack_0, ack => zeropad_same_CP_159_elements(349)); -- 
    -- CP-element group 350:  join  fork  transition  input  output  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	414 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (24) 
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_plus_offset/sum_rename_ack
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/word_access_start/$entry
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_word_addrgen/$entry
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_complete/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_word_addrgen/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_word_addrgen/root_register_ack
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_word_addrgen/root_register_req
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_complete/ack
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/word_access_start/word_0/rr
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/word_access_start/word_0/$entry
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_plus_offset/sum_rename_req
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_plus_offset/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_plus_offset/$entry
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_addr_resize/base_resize_ack
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_addr_resize/base_resize_req
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_addr_resize/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_addr_resize/$entry
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_address_resized
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_root_address_calculated
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_word_address_calculated
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_base_address_calculated
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_sample_start_
      -- 
    ack_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_957_final_reg_ack_1, ack => zeropad_same_CP_159_elements(350)); -- 
    rr_2153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(350), ack => ptr_deref_961_load_0_req_0); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351:  members (5) 
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/word_access_start/word_0/$exit
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/word_access_start/$exit
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Sample/word_access_start/word_0/ra
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_sample_completed_
      -- 
    ra_2154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_961_load_0_ack_0, ack => zeropad_same_CP_159_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	414 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: 	355 
    -- CP-element group 352: 	357 
    -- CP-element group 352: 	359 
    -- CP-element group 352: 	361 
    -- CP-element group 352: 	363 
    -- CP-element group 352: 	365 
    -- CP-element group 352: 	367 
    -- CP-element group 352:  members (33) 
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/ptr_deref_961_Merge/merge_req
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/word_access_complete/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/ptr_deref_961_Merge/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/ptr_deref_961_Merge/merge_ack
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/ptr_deref_961_Merge/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_update_completed_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/word_access_complete/word_0/ca
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/word_access_complete/word_0/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Sample/rr
      -- 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_961_load_0_ack_1, ack => zeropad_same_CP_159_elements(352)); -- 
    rr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_965_inst_req_0); -- 
    rr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_975_inst_req_0); -- 
    rr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_985_inst_req_0); -- 
    rr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_995_inst_req_0); -- 
    rr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_1005_inst_req_0); -- 
    rr_2248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_1015_inst_req_0); -- 
    rr_2262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_1025_inst_req_0); -- 
    rr_2276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(352), ack => type_cast_1035_inst_req_0); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_sample_completed_
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Sample/ra
      -- 
    ra_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_965_inst_ack_0, ack => zeropad_same_CP_159_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	414 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	389 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_update_completed_
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Update/ca
      -- 
    ca_2184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_965_inst_ack_1, ack => zeropad_same_CP_159_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	352 
    -- CP-element group 355: successors 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Sample/ra
      -- 
    ra_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_0, ack => zeropad_same_CP_159_elements(355)); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	414 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	386 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Update/ca
      -- 
    ca_2198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_1, ack => zeropad_same_CP_159_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	352 
    -- CP-element group 357: successors 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Sample/ra
      -- 
    ra_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_985_inst_ack_0, ack => zeropad_same_CP_159_elements(357)); -- 
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	414 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	383 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Update/ca
      -- 
    ca_2212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_985_inst_ack_1, ack => zeropad_same_CP_159_elements(358)); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	352 
    -- CP-element group 359: successors 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Sample/ra
      -- 
    ra_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_995_inst_ack_0, ack => zeropad_same_CP_159_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	414 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	380 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Update/ca
      -- 
    ca_2226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_995_inst_ack_1, ack => zeropad_same_CP_159_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	352 
    -- CP-element group 361: successors 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Sample/ra
      -- 
    ra_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_0, ack => zeropad_same_CP_159_elements(361)); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	414 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	377 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Update/ca
      -- 
    ca_2240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_1, ack => zeropad_same_CP_159_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	352 
    -- CP-element group 363: successors 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Sample/ra
      -- 
    ra_2249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_0, ack => zeropad_same_CP_159_elements(363)); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	414 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	374 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Update/ca
      -- 
    ca_2254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_1, ack => zeropad_same_CP_159_elements(364)); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	352 
    -- CP-element group 365: successors 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Sample/ra
      -- 
    ra_2263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_0, ack => zeropad_same_CP_159_elements(365)); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	414 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	371 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Update/ca
      -- 
    ca_2268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_1, ack => zeropad_same_CP_159_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	352 
    -- CP-element group 367: successors 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Sample/ra
      -- 
    ra_2277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_0, ack => zeropad_same_CP_159_elements(367)); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	414 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Update/ca
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Sample/req
      -- 
    ca_2282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_1, ack => zeropad_same_CP_159_elements(368)); -- 
    req_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(368), ack => WPIPE_ConvTranspose_output_pipe_1037_inst_req_0); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_update_start_
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Sample/ack
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Update/req
      -- 
    ack_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1037_inst_ack_0, ack => zeropad_same_CP_159_elements(369)); -- 
    req_2295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(369), ack => WPIPE_ConvTranspose_output_pipe_1037_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1037_Update/ack
      -- 
    ack_2296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1037_inst_ack_1, ack => zeropad_same_CP_159_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	366 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Sample/req
      -- 
    req_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(371), ack => WPIPE_ConvTranspose_output_pipe_1040_inst_req_0); -- 
    zeropad_same_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(366) & zeropad_same_CP_159_elements(370);
      gj_zeropad_same_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_update_start_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Sample/ack
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Update/req
      -- 
    ack_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1040_inst_ack_0, ack => zeropad_same_CP_159_elements(372)); -- 
    req_2309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(372), ack => WPIPE_ConvTranspose_output_pipe_1040_inst_req_1); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1040_Update/ack
      -- 
    ack_2310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1040_inst_ack_1, ack => zeropad_same_CP_159_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	364 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Sample/req
      -- 
    req_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(374), ack => WPIPE_ConvTranspose_output_pipe_1043_inst_req_0); -- 
    zeropad_same_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(364) & zeropad_same_CP_159_elements(373);
      gj_zeropad_same_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_update_start_
      -- CP-element group 375: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Sample/ack
      -- CP-element group 375: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Update/req
      -- 
    ack_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1043_inst_ack_0, ack => zeropad_same_CP_159_elements(375)); -- 
    req_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(375), ack => WPIPE_ConvTranspose_output_pipe_1043_inst_req_1); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1043_Update/ack
      -- 
    ack_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1043_inst_ack_1, ack => zeropad_same_CP_159_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	362 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Sample/req
      -- 
    req_2332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(377), ack => WPIPE_ConvTranspose_output_pipe_1046_inst_req_0); -- 
    zeropad_same_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(362) & zeropad_same_CP_159_elements(376);
      gj_zeropad_same_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_update_start_
      -- CP-element group 378: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Update/req
      -- 
    ack_2333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1046_inst_ack_0, ack => zeropad_same_CP_159_elements(378)); -- 
    req_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(378), ack => WPIPE_ConvTranspose_output_pipe_1046_inst_req_1); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1046_Update/ack
      -- 
    ack_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1046_inst_ack_1, ack => zeropad_same_CP_159_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	360 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Sample/req
      -- 
    req_2346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(380), ack => WPIPE_ConvTranspose_output_pipe_1049_inst_req_0); -- 
    zeropad_same_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(360) & zeropad_same_CP_159_elements(379);
      gj_zeropad_same_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (6) 
      -- CP-element group 381: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_update_start_
      -- CP-element group 381: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Sample/ack
      -- CP-element group 381: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Update/$entry
      -- CP-element group 381: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Update/req
      -- 
    ack_2347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1049_inst_ack_0, ack => zeropad_same_CP_159_elements(381)); -- 
    req_2351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(381), ack => WPIPE_ConvTranspose_output_pipe_1049_inst_req_1); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1049_Update/ack
      -- 
    ack_2352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1049_inst_ack_1, ack => zeropad_same_CP_159_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	358 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Sample/req
      -- 
    req_2360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(383), ack => WPIPE_ConvTranspose_output_pipe_1052_inst_req_0); -- 
    zeropad_same_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(358) & zeropad_same_CP_159_elements(382);
      gj_zeropad_same_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  transition  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_update_start_
      -- CP-element group 384: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Sample/ack
      -- CP-element group 384: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Update/req
      -- 
    ack_2361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1052_inst_ack_0, ack => zeropad_same_CP_159_elements(384)); -- 
    req_2365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(384), ack => WPIPE_ConvTranspose_output_pipe_1052_inst_req_1); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1052_Update/ack
      -- 
    ack_2366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1052_inst_ack_1, ack => zeropad_same_CP_159_elements(385)); -- 
    -- CP-element group 386:  join  transition  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	356 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_sample_start_
      -- CP-element group 386: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Sample/req
      -- 
    req_2374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(386), ack => WPIPE_ConvTranspose_output_pipe_1055_inst_req_0); -- 
    zeropad_same_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(356) & zeropad_same_CP_159_elements(385);
      gj_zeropad_same_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (6) 
      -- CP-element group 387: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_update_start_
      -- CP-element group 387: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Sample/ack
      -- CP-element group 387: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Update/req
      -- 
    ack_2375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1055_inst_ack_0, ack => zeropad_same_CP_159_elements(387)); -- 
    req_2379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(387), ack => WPIPE_ConvTranspose_output_pipe_1055_inst_req_1); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1055_Update/ack
      -- 
    ack_2380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1055_inst_ack_1, ack => zeropad_same_CP_159_elements(388)); -- 
    -- CP-element group 389:  join  transition  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	354 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Sample/req
      -- 
    req_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(389), ack => WPIPE_ConvTranspose_output_pipe_1058_inst_req_0); -- 
    zeropad_same_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(354) & zeropad_same_CP_159_elements(388);
      gj_zeropad_same_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_update_start_
      -- CP-element group 390: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Update/req
      -- 
    ack_2389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1058_inst_ack_0, ack => zeropad_same_CP_159_elements(390)); -- 
    req_2393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(390), ack => WPIPE_ConvTranspose_output_pipe_1058_inst_req_1); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/WPIPE_ConvTranspose_output_pipe_1058_Update/ack
      -- 
    ack_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1058_inst_ack_1, ack => zeropad_same_CP_159_elements(391)); -- 
    -- CP-element group 392:  branch  join  transition  place  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	347 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392: 	394 
    -- CP-element group 392:  members (10) 
      -- CP-element group 392: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071__exit__
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072__entry__
      -- CP-element group 392: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/$exit
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072_dead_link/$entry
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072_eval_test/$entry
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072_eval_test/$exit
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072_eval_test/branch_req
      -- CP-element group 392: 	 branch_block_stmt_38/R_exitcond1_1073_place
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072_if_link/$entry
      -- CP-element group 392: 	 branch_block_stmt_38/if_stmt_1072_else_link/$entry
      -- 
    branch_req_2402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(392), ack => if_stmt_1072_branch_req_0); -- 
    zeropad_same_cp_element_group_392: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_392"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(347) & zeropad_same_CP_159_elements(391);
      gj_zeropad_same_cp_element_group_392 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(392), clk => clk, reset => reset); --
    end block;
    -- CP-element group 393:  merge  transition  place  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	415 
    -- CP-element group 393:  members (13) 
      -- CP-element group 393: 	 branch_block_stmt_38/merge_stmt_1078__exit__
      -- CP-element group 393: 	 branch_block_stmt_38/forx_xend444x_xloopexit_forx_xend444
      -- CP-element group 393: 	 branch_block_stmt_38/if_stmt_1072_if_link/$exit
      -- CP-element group 393: 	 branch_block_stmt_38/if_stmt_1072_if_link/if_choice_transition
      -- CP-element group 393: 	 branch_block_stmt_38/forx_xbody371_forx_xend444x_xloopexit
      -- CP-element group 393: 	 branch_block_stmt_38/forx_xbody371_forx_xend444x_xloopexit_PhiReq/$entry
      -- CP-element group 393: 	 branch_block_stmt_38/forx_xbody371_forx_xend444x_xloopexit_PhiReq/$exit
      -- CP-element group 393: 	 branch_block_stmt_38/merge_stmt_1078_PhiReqMerge
      -- CP-element group 393: 	 branch_block_stmt_38/merge_stmt_1078_PhiAck/$entry
      -- CP-element group 393: 	 branch_block_stmt_38/merge_stmt_1078_PhiAck/$exit
      -- CP-element group 393: 	 branch_block_stmt_38/merge_stmt_1078_PhiAck/dummy
      -- CP-element group 393: 	 branch_block_stmt_38/forx_xend444x_xloopexit_forx_xend444_PhiReq/$entry
      -- CP-element group 393: 	 branch_block_stmt_38/forx_xend444x_xloopexit_forx_xend444_PhiReq/$exit
      -- 
    if_choice_transition_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1072_branch_ack_1, ack => zeropad_same_CP_159_elements(393)); -- 
    -- CP-element group 394:  fork  transition  place  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	392 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	410 
    -- CP-element group 394: 	411 
    -- CP-element group 394:  members (12) 
      -- CP-element group 394: 	 branch_block_stmt_38/if_stmt_1072_else_link/$exit
      -- CP-element group 394: 	 branch_block_stmt_38/if_stmt_1072_else_link/else_choice_transition
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Sample/rr
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1072_branch_ack_0, ack => zeropad_same_CP_159_elements(394)); -- 
    rr_2617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(394), ack => type_cast_950_inst_req_0); -- 
    cr_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(394), ack => type_cast_950_inst_req_1); -- 
    -- CP-element group 395:  merge  branch  transition  place  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	64 
    -- CP-element group 395: 	107 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	109 
    -- CP-element group 395: 	110 
    -- CP-element group 395:  members (25) 
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458_eval_test/branch_req
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_242__exit__
      -- CP-element group 395: 	 branch_block_stmt_38/forx_xcond171x_xpreheader_bbx_xnph465
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_451__exit__
      -- CP-element group 395: 	 branch_block_stmt_38/assign_stmt_457__entry__
      -- CP-element group 395: 	 branch_block_stmt_38/assign_stmt_457__exit__
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458__entry__
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458_eval_test/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458_else_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458_eval_test/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/R_cmp264448_459_place
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458_dead_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/if_stmt_458_if_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/assign_stmt_457/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/assign_stmt_457/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_242_PhiReqMerge
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_242_PhiAck/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_242_PhiAck/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_242_PhiAck/dummy
      -- CP-element group 395: 	 branch_block_stmt_38/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_451_PhiReqMerge
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_451_PhiAck/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_451_PhiAck/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/merge_stmt_451_PhiAck/dummy
      -- 
    branch_req_1018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(395), ack => if_stmt_458_branch_req_0); -- 
    zeropad_same_CP_159_elements(395) <= OrReduce(zeropad_same_CP_159_elements(64) & zeropad_same_CP_159_elements(107));
    -- CP-element group 396:  transition  output  delay-element  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	66 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	400 
    -- CP-element group 396:  members (5) 
      -- CP-element group 396: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/$exit
      -- CP-element group 396: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_282/$exit
      -- CP-element group 396: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/$exit
      -- CP-element group 396: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_286_konst_delay_trans
      -- CP-element group 396: 	 branch_block_stmt_38/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_req
      -- 
    phi_stmt_282_req_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_282_req_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(396), ack => phi_stmt_282_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(396) is a control-delay.
    cp_element_396_delay: control_delay_element  generic map(name => " 396_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(66), ack => zeropad_same_CP_159_elements(396), clk => clk, reset =>reset);
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	108 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397:  members (2) 
      -- CP-element group 397: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Sample/ra
      -- 
    ra_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_288_inst_ack_0, ack => zeropad_same_CP_159_elements(397)); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	108 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (2) 
      -- CP-element group 398: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/Update/ca
      -- 
    ca_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_288_inst_ack_1, ack => zeropad_same_CP_159_elements(398)); -- 
    -- CP-element group 399:  join  transition  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (6) 
      -- CP-element group 399: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_sources/type_cast_288/SplitProtocol/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_282/phi_stmt_282_req
      -- 
    phi_stmt_282_req_2481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_282_req_2481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(399), ack => phi_stmt_282_req_1); -- 
    zeropad_same_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(397) & zeropad_same_CP_159_elements(398);
      gj_zeropad_same_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  merge  transition  place  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	396 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_38/merge_stmt_281_PhiReqMerge
      -- CP-element group 400: 	 branch_block_stmt_38/merge_stmt_281_PhiAck/$entry
      -- 
    zeropad_same_CP_159_elements(400) <= OrReduce(zeropad_same_CP_159_elements(396) & zeropad_same_CP_159_elements(399));
    -- CP-element group 401:  fork  transition  place  input  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	67 
    -- CP-element group 401: 	68 
    -- CP-element group 401: 	70 
    -- CP-element group 401: 	71 
    -- CP-element group 401: 	74 
    -- CP-element group 401: 	78 
    -- CP-element group 401: 	82 
    -- CP-element group 401: 	86 
    -- CP-element group 401: 	90 
    -- CP-element group 401: 	94 
    -- CP-element group 401: 	98 
    -- CP-element group 401: 	102 
    -- CP-element group 401: 	105 
    -- CP-element group 401:  members (56) 
      -- CP-element group 401: 	 branch_block_stmt_38/merge_stmt_281__exit__
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444__entry__
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_resized_1
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_scaled_1
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_computed_1
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_resize_1/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_resize_1/$exit
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_resize_1/index_resize_req
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_resize_1/index_resize_ack
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_scale_1/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_scale_1/$exit
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_scale_1/scale_rename_req
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_index_scale_1/scale_rename_ack
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_update_start
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Sample/req
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/array_obj_ref_294_final_index_sum_regn_Update/req
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_complete/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/addr_of_295_complete/req
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/RPIPE_ConvTranspose_input_pipe_298_Sample/rr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_302_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_315_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_333_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_351_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_369_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_387_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_405_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/type_cast_423_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/word_access_complete/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/word_access_complete/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/assign_stmt_296_to_assign_stmt_444/ptr_deref_431_Update/word_access_complete/word_0/cr
      -- CP-element group 401: 	 branch_block_stmt_38/merge_stmt_281_PhiAck/$exit
      -- CP-element group 401: 	 branch_block_stmt_38/merge_stmt_281_PhiAck/phi_stmt_282_ack
      -- 
    phi_stmt_282_ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_282_ack_0, ack => zeropad_same_CP_159_elements(401)); -- 
    req_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => array_obj_ref_294_index_offset_req_0); -- 
    req_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => array_obj_ref_294_index_offset_req_1); -- 
    req_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => addr_of_295_final_reg_req_1); -- 
    rr_722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_0); -- 
    cr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_302_inst_req_1); -- 
    cr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_315_inst_req_1); -- 
    cr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_333_inst_req_1); -- 
    cr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_351_inst_req_1); -- 
    cr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_369_inst_req_1); -- 
    cr_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_387_inst_req_1); -- 
    cr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_405_inst_req_1); -- 
    cr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => type_cast_423_inst_req_1); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(401), ack => ptr_deref_431_store_0_req_1); -- 
    -- CP-element group 402:  transition  output  delay-element  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	112 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	406 
    -- CP-element group 402:  members (5) 
      -- CP-element group 402: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/$exit
      -- CP-element group 402: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_502/$exit
      -- CP-element group 402: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/$exit
      -- CP-element group 402: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_506_konst_delay_trans
      -- CP-element group 402: 	 branch_block_stmt_38/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_req
      -- 
    phi_stmt_502_req_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_502_req_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(402), ack => phi_stmt_502_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(402) is a control-delay.
    cp_element_402_delay: control_delay_element  generic map(name => " 402_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(112), ack => zeropad_same_CP_159_elements(402), clk => clk, reset =>reset);
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	121 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	405 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Sample/ra
      -- 
    ra_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_0, ack => zeropad_same_CP_159_elements(403)); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	121 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (2) 
      -- CP-element group 404: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/Update/ca
      -- 
    ca_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_1, ack => zeropad_same_CP_159_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	403 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (6) 
      -- CP-element group 405: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_sources/type_cast_508/SplitProtocol/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_502/phi_stmt_502_req
      -- 
    phi_stmt_502_req_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_502_req_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(405), ack => phi_stmt_502_req_1); -- 
    zeropad_same_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(403) & zeropad_same_CP_159_elements(404);
      gj_zeropad_same_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  merge  transition  place  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	402 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_38/merge_stmt_501_PhiReqMerge
      -- CP-element group 406: 	 branch_block_stmt_38/merge_stmt_501_PhiAck/$entry
      -- 
    zeropad_same_CP_159_elements(406) <= OrReduce(zeropad_same_CP_159_elements(402) & zeropad_same_CP_159_elements(405));
    -- CP-element group 407:  fork  transition  place  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	113 
    -- CP-element group 407: 	114 
    -- CP-element group 407: 	116 
    -- CP-element group 407: 	118 
    -- CP-element group 407:  members (29) 
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_complete/req
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/merge_stmt_501__exit__
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532__entry__
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_update_start_
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Update/req
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Sample/req
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_final_index_sum_regn_update_start
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_scale_1/scale_rename_ack
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_scale_1/scale_rename_req
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_scale_1/$exit
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_scale_1/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/word_access_complete/word_0/cr
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_resize_1/index_resize_ack
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_resize_1/index_resize_req
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_resize_1/$exit
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/word_access_complete/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_resize_1/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_computed_1
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_scaled_1
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/word_access_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/array_obj_ref_514_index_resized_1
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/ptr_deref_518_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/addr_of_515_update_start_
      -- CP-element group 407: 	 branch_block_stmt_38/assign_stmt_516_to_assign_stmt_532/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/merge_stmt_501_PhiAck/$exit
      -- CP-element group 407: 	 branch_block_stmt_38/merge_stmt_501_PhiAck/phi_stmt_502_ack
      -- 
    phi_stmt_502_ack_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_502_ack_0, ack => zeropad_same_CP_159_elements(407)); -- 
    req_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(407), ack => addr_of_515_final_reg_req_1); -- 
    req_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(407), ack => array_obj_ref_514_index_offset_req_1); -- 
    req_1074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(407), ack => array_obj_ref_514_index_offset_req_0); -- 
    cr_1144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(407), ack => ptr_deref_518_store_0_req_1); -- 
    -- CP-element group 408:  merge  fork  transition  place  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	110 
    -- CP-element group 408: 	120 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	122 
    -- CP-element group 408: 	123 
    -- CP-element group 408:  members (13) 
      -- CP-element group 408: 	 branch_block_stmt_38/merge_stmt_541__exit__
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544__entry__
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Update/ccr
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Update/$entry
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Sample/crr
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_update_start_
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/call_stmt_544_sample_start_
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_544/$entry
      -- CP-element group 408: 	 branch_block_stmt_38/merge_stmt_541_PhiReqMerge
      -- CP-element group 408: 	 branch_block_stmt_38/merge_stmt_541_PhiAck/$entry
      -- CP-element group 408: 	 branch_block_stmt_38/merge_stmt_541_PhiAck/$exit
      -- CP-element group 408: 	 branch_block_stmt_38/merge_stmt_541_PhiAck/dummy
      -- 
    ccr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(408), ack => call_stmt_544_call_req_1); -- 
    crr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(408), ack => call_stmt_544_call_req_0); -- 
    zeropad_same_CP_159_elements(408) <= OrReduce(zeropad_same_CP_159_elements(110) & zeropad_same_CP_159_elements(120));
    -- CP-element group 409:  transition  output  delay-element  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	346 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	413 
    -- CP-element group 409:  members (5) 
      -- CP-element group 409: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/$exit
      -- CP-element group 409: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_944/$exit
      -- CP-element group 409: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/$exit
      -- CP-element group 409: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_948_konst_delay_trans
      -- CP-element group 409: 	 branch_block_stmt_38/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_req
      -- 
    phi_stmt_944_req_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_944_req_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(409), ack => phi_stmt_944_req_0); -- 
    -- Element group zeropad_same_CP_159_elements(409) is a control-delay.
    cp_element_409_delay: control_delay_element  generic map(name => " 409_delay", delay_value => 1)  port map(req => zeropad_same_CP_159_elements(346), ack => zeropad_same_CP_159_elements(409), clk => clk, reset =>reset);
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	394 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	412 
    -- CP-element group 410:  members (2) 
      -- CP-element group 410: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Sample/ra
      -- 
    ra_2618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_950_inst_ack_0, ack => zeropad_same_CP_159_elements(410)); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	394 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (2) 
      -- CP-element group 411: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/Update/ca
      -- 
    ca_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_950_inst_ack_1, ack => zeropad_same_CP_159_elements(411)); -- 
    -- CP-element group 412:  join  transition  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	410 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/$exit
      -- CP-element group 412: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/$exit
      -- CP-element group 412: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/$exit
      -- CP-element group 412: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/$exit
      -- CP-element group 412: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_sources/type_cast_950/SplitProtocol/$exit
      -- CP-element group 412: 	 branch_block_stmt_38/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_944/phi_stmt_944_req
      -- 
    phi_stmt_944_req_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_944_req_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(412), ack => phi_stmt_944_req_1); -- 
    zeropad_same_cp_element_group_412: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_412"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_159_elements(410) & zeropad_same_CP_159_elements(411);
      gj_zeropad_same_cp_element_group_412 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_159_elements(412), clk => clk, reset => reset); --
    end block;
    -- CP-element group 413:  merge  transition  place  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	409 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (2) 
      -- CP-element group 413: 	 branch_block_stmt_38/merge_stmt_943_PhiReqMerge
      -- CP-element group 413: 	 branch_block_stmt_38/merge_stmt_943_PhiAck/$entry
      -- 
    zeropad_same_CP_159_elements(413) <= OrReduce(zeropad_same_CP_159_elements(409) & zeropad_same_CP_159_elements(412));
    -- CP-element group 414:  fork  transition  place  input  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	347 
    -- CP-element group 414: 	348 
    -- CP-element group 414: 	350 
    -- CP-element group 414: 	352 
    -- CP-element group 414: 	354 
    -- CP-element group 414: 	356 
    -- CP-element group 414: 	358 
    -- CP-element group 414: 	360 
    -- CP-element group 414: 	362 
    -- CP-element group 414: 	364 
    -- CP-element group 414: 	366 
    -- CP-element group 414: 	368 
    -- CP-element group 414:  members (53) 
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_update_start
      -- CP-element group 414: 	 branch_block_stmt_38/merge_stmt_943__exit__
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071__entry__
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_complete/req
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/word_access_complete/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/addr_of_957_complete/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_resized_1
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_scaled_1
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_computed_1
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_resize_1/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_resize_1/$exit
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_final_index_sum_regn_Update/req
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/word_access_complete/word_0/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_scale_1/scale_rename_ack
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_scale_1/scale_rename_req
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_scale_1/$exit
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_scale_1/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_resize_1/index_resize_ack
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/array_obj_ref_956_index_resize_1/index_resize_req
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/ptr_deref_961_Update/word_access_complete/word_0/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_965_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_975_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_985_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_995_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1005_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1015_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1025_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_update_start_
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/assign_stmt_958_to_assign_stmt_1071/type_cast_1035_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_38/merge_stmt_943_PhiAck/$exit
      -- CP-element group 414: 	 branch_block_stmt_38/merge_stmt_943_PhiAck/phi_stmt_944_ack
      -- 
    phi_stmt_944_ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_944_ack_0, ack => zeropad_same_CP_159_elements(414)); -- 
    req_2099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => array_obj_ref_956_index_offset_req_0); -- 
    req_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => addr_of_957_final_reg_req_1); -- 
    req_2104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => array_obj_ref_956_index_offset_req_1); -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => ptr_deref_961_load_0_req_1); -- 
    cr_2183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_965_inst_req_1); -- 
    cr_2197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_975_inst_req_1); -- 
    cr_2211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_985_inst_req_1); -- 
    cr_2225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_995_inst_req_1); -- 
    cr_2239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_1005_inst_req_1); -- 
    cr_2253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_1015_inst_req_1); -- 
    cr_2267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_1025_inst_req_1); -- 
    cr_2281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_159_elements(414), ack => type_cast_1035_inst_req_1); -- 
    -- CP-element group 415:  merge  transition  place  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	344 
    -- CP-element group 415: 	393 
    -- CP-element group 415: successors 
    -- CP-element group 415:  members (16) 
      -- CP-element group 415: 	 $exit
      -- CP-element group 415: 	 branch_block_stmt_38/$exit
      -- CP-element group 415: 	 branch_block_stmt_38/branch_block_stmt_38__exit__
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1080__exit__
      -- CP-element group 415: 	 branch_block_stmt_38/return__
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1082__exit__
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1080_PhiReqMerge
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1080_PhiAck/$entry
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1080_PhiAck/$exit
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1080_PhiAck/dummy
      -- CP-element group 415: 	 branch_block_stmt_38/return___PhiReq/$entry
      -- CP-element group 415: 	 branch_block_stmt_38/return___PhiReq/$exit
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1082_PhiReqMerge
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1082_PhiAck/$entry
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1082_PhiAck/$exit
      -- CP-element group 415: 	 branch_block_stmt_38/merge_stmt_1082_PhiAck/dummy
      -- 
    zeropad_same_CP_159_elements(415) <= OrReduce(zeropad_same_CP_159_elements(344) & zeropad_same_CP_159_elements(393));
    zeropad_same_do_while_stmt_575_terminator_1760: loop_terminator -- 
      generic map (name => " zeropad_same_do_while_stmt_575_terminator_1760", max_iterations_in_flight =>15) 
      port map(loop_body_exit => zeropad_same_CP_159_elements(128),loop_continue => zeropad_same_CP_159_elements(295),loop_terminate => zeropad_same_CP_159_elements(294),loop_back => zeropad_same_CP_159_elements(126),loop_exit => zeropad_same_CP_159_elements(125),clk => clk, reset => reset); -- 
    phi_stmt_577_phi_seq_1248_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_159_elements(143);
      zeropad_same_CP_159_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_159_elements(146);
      zeropad_same_CP_159_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_159_elements(148);
      zeropad_same_CP_159_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_159_elements(141);
      zeropad_same_CP_159_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_159_elements(152);
      zeropad_same_CP_159_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_159_elements(153);
      zeropad_same_CP_159_elements(142) <= phi_mux_reqs(1);
      phi_stmt_577_phi_seq_1248 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_577_phi_seq_1248") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_159_elements(133), 
          phi_sample_ack => zeropad_same_CP_159_elements(139), 
          phi_update_req => zeropad_same_CP_159_elements(135), 
          phi_update_ack => zeropad_same_CP_159_elements(140), 
          phi_mux_ack => zeropad_same_CP_159_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_581_phi_seq_1292_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_159_elements(162);
      zeropad_same_CP_159_elements(165)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_159_elements(165);
      zeropad_same_CP_159_elements(166)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_159_elements(167);
      zeropad_same_CP_159_elements(163) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_159_elements(160);
      zeropad_same_CP_159_elements(169)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_159_elements(171);
      zeropad_same_CP_159_elements(170)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_159_elements(172);
      zeropad_same_CP_159_elements(161) <= phi_mux_reqs(1);
      phi_stmt_581_phi_seq_1292 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_581_phi_seq_1292") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_159_elements(156), 
          phi_sample_ack => zeropad_same_CP_159_elements(157), 
          phi_update_req => zeropad_same_CP_159_elements(158), 
          phi_update_ack => zeropad_same_CP_159_elements(159), 
          phi_mux_ack => zeropad_same_CP_159_elements(164), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_585_phi_seq_1336_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_159_elements(181);
      zeropad_same_CP_159_elements(184)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_159_elements(184);
      zeropad_same_CP_159_elements(185)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_159_elements(186);
      zeropad_same_CP_159_elements(182) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_159_elements(179);
      zeropad_same_CP_159_elements(188)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_159_elements(190);
      zeropad_same_CP_159_elements(189)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_159_elements(191);
      zeropad_same_CP_159_elements(180) <= phi_mux_reqs(1);
      phi_stmt_585_phi_seq_1336 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_585_phi_seq_1336") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_159_elements(175), 
          phi_sample_ack => zeropad_same_CP_159_elements(176), 
          phi_update_req => zeropad_same_CP_159_elements(177), 
          phi_update_ack => zeropad_same_CP_159_elements(178), 
          phi_mux_ack => zeropad_same_CP_159_elements(183), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_589_phi_seq_1390_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_159_elements(200);
      zeropad_same_CP_159_elements(203)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_159_elements(205);
      zeropad_same_CP_159_elements(204)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_159_elements(206);
      zeropad_same_CP_159_elements(201) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_159_elements(198);
      zeropad_same_CP_159_elements(207)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_159_elements(209);
      zeropad_same_CP_159_elements(208)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_159_elements(210);
      zeropad_same_CP_159_elements(199) <= phi_mux_reqs(1);
      phi_stmt_589_phi_seq_1390 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_589_phi_seq_1390") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_159_elements(194), 
          phi_sample_ack => zeropad_same_CP_159_elements(195), 
          phi_update_req => zeropad_same_CP_159_elements(196), 
          phi_update_ack => zeropad_same_CP_159_elements(197), 
          phi_mux_ack => zeropad_same_CP_159_elements(202), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_593_phi_seq_1444_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_159_elements(219);
      zeropad_same_CP_159_elements(222)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_159_elements(224);
      zeropad_same_CP_159_elements(223)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_159_elements(225);
      zeropad_same_CP_159_elements(220) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_159_elements(217);
      zeropad_same_CP_159_elements(226)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_159_elements(228);
      zeropad_same_CP_159_elements(227)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_159_elements(229);
      zeropad_same_CP_159_elements(218) <= phi_mux_reqs(1);
      phi_stmt_593_phi_seq_1444 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_593_phi_seq_1444") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_159_elements(213), 
          phi_sample_ack => zeropad_same_CP_159_elements(214), 
          phi_update_req => zeropad_same_CP_159_elements(215), 
          phi_update_ack => zeropad_same_CP_159_elements(216), 
          phi_mux_ack => zeropad_same_CP_159_elements(221), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_597_phi_seq_1488_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_159_elements(238);
      zeropad_same_CP_159_elements(241)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_159_elements(241);
      zeropad_same_CP_159_elements(242)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_159_elements(243);
      zeropad_same_CP_159_elements(239) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_159_elements(236);
      zeropad_same_CP_159_elements(245)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_159_elements(247);
      zeropad_same_CP_159_elements(246)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_159_elements(248);
      zeropad_same_CP_159_elements(237) <= phi_mux_reqs(1);
      phi_stmt_597_phi_seq_1488 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_597_phi_seq_1488") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_159_elements(232), 
          phi_sample_ack => zeropad_same_CP_159_elements(233), 
          phi_update_req => zeropad_same_CP_159_elements(234), 
          phi_update_ack => zeropad_same_CP_159_elements(235), 
          phi_mux_ack => zeropad_same_CP_159_elements(240), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1200_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= zeropad_same_CP_159_elements(129);
        preds(1)  <= zeropad_same_CP_159_elements(130);
        entry_tmerge_1200 : transition_merge -- 
          generic map(name => " entry_tmerge_1200")
          port map (preds => preds, symbol_out => zeropad_same_CP_159_elements(131));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_725_wire : std_logic_vector(15 downto 0);
    signal MUX_747_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_679_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_721_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_743_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_770_wire : std_logic_vector(0 downto 0);
    signal R_indvar469_513_resized : std_logic_vector(13 downto 0);
    signal R_indvar469_513_scaled : std_logic_vector(13 downto 0);
    signal R_indvar489_293_resized : std_logic_vector(13 downto 0);
    signal R_indvar489_293_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_955_resized : std_logic_vector(13 downto 0);
    signal R_indvar_955_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_561_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_665_665_delayed_1_0_671 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_749_749_delayed_1_0_761 : std_logic_vector(15 downto 0);
    signal add131_321 : std_logic_vector(63 downto 0);
    signal add137_339 : std_logic_vector(63 downto 0);
    signal add143_357 : std_logic_vector(63 downto 0);
    signal add149_375 : std_logic_vector(63 downto 0);
    signal add155_393 : std_logic_vector(63 downto 0);
    signal add161_411 : std_logic_vector(63 downto 0);
    signal add167_429 : std_logic_vector(63 downto 0);
    signal add_dest_dim0_589 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_567 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_567_591_buffered : std_logic_vector(15 downto 0);
    signal add_dest_dim1_593 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_570 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_570_595_buffered : std_logic_vector(15 downto 0);
    signal add_out_626 : std_logic_vector(15 downto 0);
    signal add_src_597 : std_logic_vector(31 downto 0);
    signal add_src_init_574 : std_logic_vector(31 downto 0);
    signal array_obj_ref_294_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_294_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_294_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_294_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_294_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_294_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_514_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_514_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_514_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_514_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_514_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_514_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_632_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_632_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_632_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_632_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_632_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_632_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_644_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_644_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_644_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_644_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_644_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_644_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_956_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_956_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_956_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_956_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_956_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_956_root_address : std_logic_vector(13 downto 0);
    signal arrayidx269_516 : std_logic_vector(31 downto 0);
    signal arrayidx376_958 : std_logic_vector(31 downto 0);
    signal arrayidx_296 : std_logic_vector(31 downto 0);
    signal call10_80 : std_logic_vector(7 downto 0);
    signal call110_117 : std_logic_vector(7 downto 0);
    signal call1124_155 : std_logic_vector(7 downto 0);
    signal call1128_167 : std_logic_vector(7 downto 0);
    signal call115_130 : std_logic_vector(7 downto 0);
    signal call119_142 : std_logic_vector(7 downto 0);
    signal call124_299 : std_logic_vector(7 downto 0);
    signal call128_312 : std_logic_vector(7 downto 0);
    signal call133_180 : std_logic_vector(7 downto 0);
    signal call134_330 : std_logic_vector(7 downto 0);
    signal call140_348 : std_logic_vector(7 downto 0);
    signal call146_366 : std_logic_vector(7 downto 0);
    signal call14_92 : std_logic_vector(7 downto 0);
    signal call152_384 : std_logic_vector(7 downto 0);
    signal call158_402 : std_logic_vector(7 downto 0);
    signal call164_420 : std_logic_vector(7 downto 0);
    signal call19_105 : std_logic_vector(7 downto 0);
    signal call233_544 : std_logic_vector(63 downto 0);
    signal call297_777 : std_logic_vector(63 downto 0);
    signal call2_55 : std_logic_vector(7 downto 0);
    signal call5_67 : std_logic_vector(7 downto 0);
    signal call_41 : std_logic_vector(7 downto 0);
    signal cmp264448_457 : std_logic_vector(0 downto 0);
    signal cmp264449_899 : std_logic_vector(0 downto 0);
    signal cmp467_233 : std_logic_vector(0 downto 0);
    signal cmp_dim0_682 : std_logic_vector(0 downto 0);
    signal cmp_dim1_676 : std_logic_vector(0 downto 0);
    signal cmp_dim2_666 : std_logic_vector(0 downto 0);
    signal continue_flag_772 : std_logic_vector(0 downto 0);
    signal conv1125_159 : std_logic_vector(15 downto 0);
    signal conv113_121 : std_logic_vector(15 downto 0);
    signal conv116_134 : std_logic_vector(15 downto 0);
    signal conv11_84 : std_logic_vector(15 downto 0);
    signal conv122_146 : std_logic_vector(15 downto 0);
    signal conv125_303 : std_logic_vector(63 downto 0);
    signal conv130_316 : std_logic_vector(63 downto 0);
    signal conv131_171 : std_logic_vector(15 downto 0);
    signal conv134_184 : std_logic_vector(15 downto 0);
    signal conv136_334 : std_logic_vector(63 downto 0);
    signal conv142_352 : std_logic_vector(63 downto 0);
    signal conv148_370 : std_logic_vector(63 downto 0);
    signal conv154_388 : std_logic_vector(63 downto 0);
    signal conv160_406 : std_logic_vector(63 downto 0);
    signal conv166_424 : std_logic_vector(63 downto 0);
    signal conv17_96 : std_logic_vector(15 downto 0);
    signal conv1_46 : std_logic_vector(15 downto 0);
    signal conv20_109 : std_logic_vector(15 downto 0);
    signal conv276_783 : std_logic_vector(63 downto 0);
    signal conv298_788 : std_logic_vector(63 downto 0);
    signal conv305_798 : std_logic_vector(7 downto 0);
    signal conv311_808 : std_logic_vector(7 downto 0);
    signal conv317_818 : std_logic_vector(7 downto 0);
    signal conv323_828 : std_logic_vector(7 downto 0);
    signal conv329_838 : std_logic_vector(7 downto 0);
    signal conv335_848 : std_logic_vector(7 downto 0);
    signal conv341_858 : std_logic_vector(7 downto 0);
    signal conv347_868 : std_logic_vector(7 downto 0);
    signal conv381_966 : std_logic_vector(7 downto 0);
    signal conv387_976 : std_logic_vector(7 downto 0);
    signal conv393_986 : std_logic_vector(7 downto 0);
    signal conv399_996 : std_logic_vector(7 downto 0);
    signal conv3_59 : std_logic_vector(15 downto 0);
    signal conv405_1006 : std_logic_vector(7 downto 0);
    signal conv411_1016 : std_logic_vector(7 downto 0);
    signal conv417_1026 : std_logic_vector(7 downto 0);
    signal conv423_1036 : std_logic_vector(7 downto 0);
    signal conv8_71 : std_logic_vector(15 downto 0);
    signal dim0_end_766 : std_logic_vector(0 downto 0);
    signal dim2_limit_658 : std_logic_vector(15 downto 0);
    signal dim2_limit_658_delayed_1_0_661 : std_logic_vector(15 downto 0);
    signal exitcond1_1071 : std_logic_vector(0 downto 0);
    signal exitcond2_444 : std_logic_vector(0 downto 0);
    signal exitcond_532 : std_logic_vector(0 downto 0);
    signal i1_638 : std_logic_vector(63 downto 0);
    signal iNsTr_111_928 : std_logic_vector(63 downto 0);
    signal iNsTr_19_266 : std_logic_vector(63 downto 0);
    signal iNsTr_52_486 : std_logic_vector(63 downto 0);
    signal indvar469_502 : std_logic_vector(63 downto 0);
    signal indvar489_282 : std_logic_vector(63 downto 0);
    signal indvar_944 : std_logic_vector(63 downto 0);
    signal indvarx_xnext470_527 : std_logic_vector(63 downto 0);
    signal indvarx_xnext490_439 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1066 : std_logic_vector(63 downto 0);
    signal inp_d0_64 : std_logic_vector(15 downto 0);
    signal inp_d1_89 : std_logic_vector(15 downto 0);
    signal inp_d232_194 : std_logic_vector(31 downto 0);
    signal inp_d2_114 : std_logic_vector(15 downto 0);
    signal input_dim0_577 : std_logic_vector(15 downto 0);
    signal input_dim0_init_549 : std_logic_vector(15 downto 0);
    signal input_dim1_581 : std_logic_vector(15 downto 0);
    signal input_dim1_init_553 : std_logic_vector(15 downto 0);
    signal input_dim2_585 : std_logic_vector(15 downto 0);
    signal input_dim2_init_557 : std_logic_vector(15 downto 0);
    signal input_int1_203 : std_logic_vector(31 downto 0);
    signal input_int_199 : std_logic_vector(15 downto 0);
    signal input_size_208 : std_logic_vector(31 downto 0);
    signal iv1_634 : std_logic_vector(31 downto 0);
    signal konst_562_wire_constant : std_logic_vector(15 downto 0);
    signal konst_624_wire_constant : std_logic_vector(15 downto 0);
    signal konst_656_wire_constant : std_logic_vector(15 downto 0);
    signal konst_669_wire_constant : std_logic_vector(15 downto 0);
    signal konst_685_wire_constant : std_logic_vector(15 downto 0);
    signal konst_690_wire_constant : std_logic_vector(15 downto 0);
    signal konst_695_wire_constant : std_logic_vector(15 downto 0);
    signal konst_700_wire_constant : std_logic_vector(15 downto 0);
    signal konst_705_wire_constant : std_logic_vector(15 downto 0);
    signal konst_713_wire_constant : std_logic_vector(31 downto 0);
    signal konst_738_wire_constant : std_logic_vector(15 downto 0);
    signal konst_759_wire_constant : std_logic_vector(15 downto 0);
    signal nao1_611 : std_logic_vector(15 downto 0);
    signal nao2_616 : std_logic_vector(15 downto 0);
    signal nao3_621 : std_logic_vector(15 downto 0);
    signal nao_606 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_734 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_734_592_buffered : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_728 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_728_596_buffered : std_logic_vector(15 downto 0);
    signal next_add_src_715 : std_logic_vector(31 downto 0);
    signal next_add_src_715_600_buffered : std_logic_vector(31 downto 0);
    signal next_input_dim0_756 : std_logic_vector(15 downto 0);
    signal next_input_dim0_756_580_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim1_750 : std_logic_vector(15 downto 0);
    signal next_input_dim1_750_584_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim2_740 : std_logic_vector(15 downto 0);
    signal next_input_dim2_740_588_buffered : std_logic_vector(15 downto 0);
    signal nid1_true1_707 : std_logic_vector(15 downto 0);
    signal nid1_true4_710 : std_logic_vector(15 downto 0);
    signal nid1_true4_711_delayed_1_0_718 : std_logic_vector(15 downto 0);
    signal nid1_true_702 : std_logic_vector(15 downto 0);
    signal nid2_false1_697 : std_logic_vector(15 downto 0);
    signal nid2_false_692 : std_logic_vector(15 downto 0);
    signal nid2_true_687 : std_logic_vector(15 downto 0);
    signal out_d0_139 : std_logic_vector(15 downto 0);
    signal out_d1_164 : std_logic_vector(15 downto 0);
    signal out_d232_212 : std_logic_vector(31 downto 0);
    signal out_d2_189 : std_logic_vector(15 downto 0);
    signal out_int1_221 : std_logic_vector(31 downto 0);
    signal out_int_217 : std_logic_vector(15 downto 0);
    signal output_size_226 : std_logic_vector(31 downto 0);
    signal ov_646 : std_logic_vector(31 downto 0);
    signal ov_647_delayed_6_0_649 : std_logic_vector(31 downto 0);
    signal pad_564 : std_logic_vector(15 downto 0);
    signal ptr_deref_431_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_431_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_431_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_431_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_431_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_431_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_518_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_518_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_518_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_518_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_518_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_518_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_637_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_637_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_637_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_637_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_637_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_651_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_651_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_651_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_651_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_651_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_651_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_961_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_961_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_961_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_961_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_961_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl114_127 : std_logic_vector(15 downto 0);
    signal shl123_152 : std_logic_vector(15 downto 0);
    signal shl127_309 : std_logic_vector(63 downto 0);
    signal shl132_177 : std_logic_vector(15 downto 0);
    signal shl133_327 : std_logic_vector(63 downto 0);
    signal shl139_345 : std_logic_vector(63 downto 0);
    signal shl145_363 : std_logic_vector(63 downto 0);
    signal shl151_381 : std_logic_vector(63 downto 0);
    signal shl157_399 : std_logic_vector(63 downto 0);
    signal shl163_417 : std_logic_vector(63 downto 0);
    signal shl18_102 : std_logic_vector(15 downto 0);
    signal shl9_77 : std_logic_vector(15 downto 0);
    signal shl_52 : std_logic_vector(15 downto 0);
    signal shr308_804 : std_logic_vector(63 downto 0);
    signal shr314_814 : std_logic_vector(63 downto 0);
    signal shr320_824 : std_logic_vector(63 downto 0);
    signal shr326_834 : std_logic_vector(63 downto 0);
    signal shr332_844 : std_logic_vector(63 downto 0);
    signal shr338_854 : std_logic_vector(63 downto 0);
    signal shr344_864 : std_logic_vector(63 downto 0);
    signal shr384_972 : std_logic_vector(63 downto 0);
    signal shr390_982 : std_logic_vector(63 downto 0);
    signal shr396_992 : std_logic_vector(63 downto 0);
    signal shr402_1002 : std_logic_vector(63 downto 0);
    signal shr408_1012 : std_logic_vector(63 downto 0);
    signal shr414_1022 : std_logic_vector(63 downto 0);
    signal shr420_1032 : std_logic_vector(63 downto 0);
    signal sub_793 : std_logic_vector(63 downto 0);
    signal tmp377_962 : std_logic_vector(63 downto 0);
    signal tmp464_912 : std_logic_vector(31 downto 0);
    signal tmp464x_xop_924 : std_logic_vector(31 downto 0);
    signal tmp465_918 : std_logic_vector(0 downto 0);
    signal tmp468_941 : std_logic_vector(63 downto 0);
    signal tmp476_470 : std_logic_vector(31 downto 0);
    signal tmp476x_xop_482 : std_logic_vector(31 downto 0);
    signal tmp477_476 : std_logic_vector(0 downto 0);
    signal tmp481_499 : std_logic_vector(63 downto 0);
    signal tmp495_250 : std_logic_vector(31 downto 0);
    signal tmp495x_xop_262 : std_logic_vector(31 downto 0);
    signal tmp496_256 : std_logic_vector(0 downto 0);
    signal tmp500_279 : std_logic_vector(63 downto 0);
    signal type_cast_1000_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_100_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1020_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_125_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_150_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_175_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_230_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_248_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_254_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_260_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_270_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_277_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_286_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_288_wire : std_logic_vector(63 downto 0);
    signal type_cast_307_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_343_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_361_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_379_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_397_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_415_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_437_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_455_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_468_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_480_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_490_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_497_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_506_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_508_wire : std_logic_vector(63 downto 0);
    signal type_cast_50_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_525_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_631_resized : std_logic_vector(13 downto 0);
    signal type_cast_631_scaled : std_logic_vector(13 downto 0);
    signal type_cast_631_wire : std_logic_vector(63 downto 0);
    signal type_cast_643_resized : std_logic_vector(13 downto 0);
    signal type_cast_643_scaled : std_logic_vector(13 downto 0);
    signal type_cast_643_wire : std_logic_vector(63 downto 0);
    signal type_cast_75_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_781_wire : std_logic_vector(63 downto 0);
    signal type_cast_786_wire : std_logic_vector(63 downto 0);
    signal type_cast_802_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_812_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_822_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_832_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_842_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_852_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_862_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_910_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_922_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_932_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_939_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_950_wire : std_logic_vector(63 downto 0);
    signal type_cast_970_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_980_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_990_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop503_272 : std_logic_vector(63 downto 0);
    signal xx_xop513_492 : std_logic_vector(63 downto 0);
    signal xx_xop_934 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    add_src_init_574 <= "00000000000000000000000000000000";
    array_obj_ref_294_constant_part_of_offset <= "00000000000000";
    array_obj_ref_294_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_294_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_294_resized_base_address <= "00000000000000";
    array_obj_ref_514_constant_part_of_offset <= "00000000000000";
    array_obj_ref_514_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_514_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_514_resized_base_address <= "00000000000000";
    array_obj_ref_632_constant_part_of_offset <= "00000000000000";
    array_obj_ref_632_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_632_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_632_resized_base_address <= "00000000000000";
    array_obj_ref_644_constant_part_of_offset <= "00000000000000";
    array_obj_ref_644_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_644_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_644_resized_base_address <= "00000000000000";
    array_obj_ref_956_constant_part_of_offset <= "00000000000000";
    array_obj_ref_956_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_956_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_956_resized_base_address <= "00000000000000";
    input_dim0_init_549 <= "0000000000000000";
    input_dim1_init_553 <= "0000000000000000";
    input_dim2_init_557 <= "0000000000000000";
    konst_562_wire_constant <= "0000000000000001";
    konst_624_wire_constant <= "0000000000000011";
    konst_656_wire_constant <= "0000000000001000";
    konst_669_wire_constant <= "0000000000000001";
    konst_685_wire_constant <= "0000000000001000";
    konst_690_wire_constant <= "0000000000000001";
    konst_695_wire_constant <= "0000000000000001";
    konst_700_wire_constant <= "0000000000000001";
    konst_705_wire_constant <= "0000000000000001";
    konst_713_wire_constant <= "00000000000000000000000000000001";
    konst_738_wire_constant <= "0000000000000000";
    konst_759_wire_constant <= "0000000000000001";
    ptr_deref_431_word_offset_0 <= "00000000000000";
    ptr_deref_518_word_offset_0 <= "00000000000000";
    ptr_deref_637_word_offset_0 <= "00000000000000";
    ptr_deref_651_word_offset_0 <= "00000000000000";
    ptr_deref_961_word_offset_0 <= "00000000000000";
    type_cast_1000_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_100_wire_constant <= "0000000000001000";
    type_cast_1010_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1020_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1064_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_125_wire_constant <= "0000000000001000";
    type_cast_150_wire_constant <= "0000000000001000";
    type_cast_175_wire_constant <= "0000000000001000";
    type_cast_230_wire_constant <= "00000000000000000000000000000111";
    type_cast_248_wire_constant <= "00000000000000000000000000000011";
    type_cast_254_wire_constant <= "00000000000000000000000000000001";
    type_cast_260_wire_constant <= "11111111111111111111111111111111";
    type_cast_270_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_286_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_307_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_325_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_343_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_361_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_379_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_397_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_415_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_455_wire_constant <= "00000000000000000000000000000011";
    type_cast_468_wire_constant <= "00000000000000000000000000000011";
    type_cast_474_wire_constant <= "00000000000000000000000000000001";
    type_cast_480_wire_constant <= "11111111111111111111111111111111";
    type_cast_490_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_497_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_506_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_50_wire_constant <= "0000000000001000";
    type_cast_520_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_525_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_75_wire_constant <= "0000000000001000";
    type_cast_802_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_812_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_822_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_832_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_842_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_852_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_862_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_897_wire_constant <= "00000000000000000000000000000111";
    type_cast_910_wire_constant <= "00000000000000000000000000000011";
    type_cast_916_wire_constant <= "00000000000000000000000000000001";
    type_cast_922_wire_constant <= "11111111111111111111111111111111";
    type_cast_932_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_939_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_948_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_970_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_980_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_990_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    phi_stmt_282: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_286_wire_constant & type_cast_288_wire;
      req <= phi_stmt_282_req_0 & phi_stmt_282_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_282",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_282_ack_0,
          idata => idata,
          odata => indvar489_282,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_282
    phi_stmt_502: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_506_wire_constant & type_cast_508_wire;
      req <= phi_stmt_502_req_0 & phi_stmt_502_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_502",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_502_ack_0,
          idata => idata,
          odata => indvar469_502,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_502
    phi_stmt_577: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim0_init_549 & next_input_dim0_756_580_buffered;
      req <= phi_stmt_577_req_0 & phi_stmt_577_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_577",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_577_ack_0,
          idata => idata,
          odata => input_dim0_577,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_577
    phi_stmt_581: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim1_init_553 & next_input_dim1_750_584_buffered;
      req <= phi_stmt_581_req_0 & phi_stmt_581_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_581",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_581_ack_0,
          idata => idata,
          odata => input_dim1_581,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_581
    phi_stmt_585: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim2_init_557 & next_input_dim2_740_588_buffered;
      req <= phi_stmt_585_req_0 & phi_stmt_585_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_585",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_585_ack_0,
          idata => idata,
          odata => input_dim2_585,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_585
    phi_stmt_589: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim0_init_567_591_buffered & next_add_dest_dim0_734_592_buffered;
      req <= phi_stmt_589_req_0 & phi_stmt_589_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_589",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_589_ack_0,
          idata => idata,
          odata => add_dest_dim0_589,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_589
    phi_stmt_593: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim1_init_570_595_buffered & next_add_dest_dim1_728_596_buffered;
      req <= phi_stmt_593_req_0 & phi_stmt_593_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_593",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_593_ack_0,
          idata => idata,
          odata => add_dest_dim1_593,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_593
    phi_stmt_597: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_src_init_574 & next_add_src_715_600_buffered;
      req <= phi_stmt_597_req_0 & phi_stmt_597_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_597",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_597_ack_0,
          idata => idata,
          odata => add_src_597,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_597
    phi_stmt_944: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_948_wire_constant & type_cast_950_wire;
      req <= phi_stmt_944_req_0 & phi_stmt_944_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_944",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_944_ack_0,
          idata => idata,
          odata => indvar_944,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_944
    -- flow-through select operator MUX_278_inst
    tmp500_279 <= xx_xop503_272 when (tmp496_256(0) /=  '0') else type_cast_277_wire_constant;
    -- flow-through select operator MUX_498_inst
    tmp481_499 <= xx_xop513_492 when (tmp477_476(0) /=  '0') else type_cast_497_wire_constant;
    -- flow-through select operator MUX_725_inst
    MUX_725_wire <= nid1_true4_711_delayed_1_0_718 when (cmp_dim1_676(0) /=  '0') else nid2_false1_697;
    -- flow-through select operator MUX_727_inst
    next_add_dest_dim1_728 <= MUX_725_wire when (NOT_u1_u1_721_wire(0) /=  '0') else add_dest_dim1_593;
    -- flow-through select operator MUX_733_inst
    next_add_dest_dim0_734 <= nid1_true1_707 when (cmp_dim0_682(0) /=  '0') else add_dest_dim0_589;
    -- flow-through select operator MUX_739_inst
    next_input_dim2_740 <= nid2_true_687 when (cmp_dim2_666(0) /=  '0') else konst_738_wire_constant;
    -- flow-through select operator MUX_747_inst
    MUX_747_wire <= pad_564 when (cmp_dim1_676(0) /=  '0') else nid2_false_692;
    -- flow-through select operator MUX_749_inst
    next_input_dim1_750 <= MUX_747_wire when (NOT_u1_u1_743_wire(0) /=  '0') else input_dim1_581;
    -- flow-through select operator MUX_755_inst
    next_input_dim0_756 <= nid1_true_702 when (cmp_dim0_682(0) /=  '0') else input_dim0_577;
    -- flow-through select operator MUX_940_inst
    tmp468_941 <= xx_xop_934 when (tmp465_918(0) /=  '0') else type_cast_939_wire_constant;
    -- interlock W_add_dest_dim0_init_565_inst
    process(pad_564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := pad_564(15 downto 0);
      add_dest_dim0_init_567 <= tmp_var; -- 
    end process;
    -- interlock W_add_dest_dim1_init_568_inst
    process(pad_564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := pad_564(15 downto 0);
      add_dest_dim1_init_570 <= tmp_var; -- 
    end process;
    W_dim2_limit_658_delayed_1_0_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dim2_limit_658_delayed_1_0_659_inst_req_0;
      W_dim2_limit_658_delayed_1_0_659_inst_ack_0<= wack(0);
      rreq(0) <= W_dim2_limit_658_delayed_1_0_659_inst_req_1;
      W_dim2_limit_658_delayed_1_0_659_inst_ack_1<= rack(0);
      W_dim2_limit_658_delayed_1_0_659_inst : InterlockBuffer generic map ( -- 
        name => "W_dim2_limit_658_delayed_1_0_659_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dim2_limit_658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dim2_limit_658_delayed_1_0_661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nid1_true4_708_inst
    process(pad_564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := pad_564(15 downto 0);
      nid1_true4_710 <= tmp_var; -- 
    end process;
    W_nid1_true4_711_delayed_1_0_716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_nid1_true4_711_delayed_1_0_716_inst_req_0;
      W_nid1_true4_711_delayed_1_0_716_inst_ack_0<= wack(0);
      rreq(0) <= W_nid1_true4_711_delayed_1_0_716_inst_req_1;
      W_nid1_true4_711_delayed_1_0_716_inst_ack_1<= rack(0);
      W_nid1_true4_711_delayed_1_0_716_inst : InterlockBuffer generic map ( -- 
        name => "W_nid1_true4_711_delayed_1_0_716_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nid1_true4_710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nid1_true4_711_delayed_1_0_718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ov_647_delayed_6_0_647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ov_647_delayed_6_0_647_inst_req_0;
      W_ov_647_delayed_6_0_647_inst_ack_0<= wack(0);
      rreq(0) <= W_ov_647_delayed_6_0_647_inst_req_1;
      W_ov_647_delayed_6_0_647_inst_ack_1<= rack(0);
      W_ov_647_delayed_6_0_647_inst : InterlockBuffer generic map ( -- 
        name => "W_ov_647_delayed_6_0_647_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ov_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ov_647_delayed_6_0_649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim0_init_567_591_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim0_init_567_591_buf_req_0;
      add_dest_dim0_init_567_591_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim0_init_567_591_buf_req_1;
      add_dest_dim0_init_567_591_buf_ack_1<= rack(0);
      add_dest_dim0_init_567_591_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim0_init_567_591_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0_init_567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim0_init_567_591_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim1_init_570_595_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim1_init_570_595_buf_req_0;
      add_dest_dim1_init_570_595_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim1_init_570_595_buf_req_1;
      add_dest_dim1_init_570_595_buf_ack_1<= rack(0);
      add_dest_dim1_init_570_595_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim1_init_570_595_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1_init_570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1_init_570_595_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_295_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_295_final_reg_req_0;
      addr_of_295_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_295_final_reg_req_1;
      addr_of_295_final_reg_ack_1<= rack(0);
      addr_of_295_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_295_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_294_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_515_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_515_final_reg_req_0;
      addr_of_515_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_515_final_reg_req_1;
      addr_of_515_final_reg_ack_1<= rack(0);
      addr_of_515_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_515_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_514_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_633_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_633_final_reg_req_0;
      addr_of_633_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_633_final_reg_req_1;
      addr_of_633_final_reg_ack_1<= rack(0);
      addr_of_633_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_633_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_632_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iv1_634,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_645_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_645_final_reg_req_0;
      addr_of_645_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_645_final_reg_req_1;
      addr_of_645_final_reg_ack_1<= rack(0);
      addr_of_645_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_645_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_644_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ov_646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_957_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_957_final_reg_req_0;
      addr_of_957_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_957_final_reg_req_1;
      addr_of_957_final_reg_ack_1<= rack(0);
      addr_of_957_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_957_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_956_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx376_958,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim0_734_592_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim0_734_592_buf_req_0;
      next_add_dest_dim0_734_592_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim0_734_592_buf_req_1;
      next_add_dest_dim0_734_592_buf_ack_1<= rack(0);
      next_add_dest_dim0_734_592_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim0_734_592_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim0_734,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim0_734_592_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim1_728_596_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim1_728_596_buf_req_0;
      next_add_dest_dim1_728_596_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim1_728_596_buf_req_1;
      next_add_dest_dim1_728_596_buf_ack_1<= rack(0);
      next_add_dest_dim1_728_596_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim1_728_596_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim1_728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim1_728_596_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_src_715_600_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_src_715_600_buf_req_0;
      next_add_src_715_600_buf_ack_0<= wack(0);
      rreq(0) <= next_add_src_715_600_buf_req_1;
      next_add_src_715_600_buf_ack_1<= rack(0);
      next_add_src_715_600_buf : InterlockBuffer generic map ( -- 
        name => "next_add_src_715_600_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_src_715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_src_715_600_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim0_756_580_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim0_756_580_buf_req_0;
      next_input_dim0_756_580_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim0_756_580_buf_req_1;
      next_input_dim0_756_580_buf_ack_1<= rack(0);
      next_input_dim0_756_580_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim0_756_580_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim0_756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim0_756_580_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim1_750_584_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim1_750_584_buf_req_0;
      next_input_dim1_750_584_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim1_750_584_buf_req_1;
      next_input_dim1_750_584_buf_ack_1<= rack(0);
      next_input_dim1_750_584_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim1_750_584_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim1_750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim1_750_584_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim2_740_588_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim2_740_588_buf_req_0;
      next_input_dim2_740_588_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim2_740_588_buf_req_1;
      next_input_dim2_740_588_buf_ack_1<= rack(0);
      next_input_dim2_740_588_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim2_740_588_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim2_740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim2_740_588_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1005_inst_req_0;
      type_cast_1005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1005_inst_req_1;
      type_cast_1005_inst_ack_1<= rack(0);
      type_cast_1005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr402_1002,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv405_1006,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1015_inst_req_0;
      type_cast_1015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1015_inst_req_1;
      type_cast_1015_inst_ack_1<= rack(0);
      type_cast_1015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr408_1012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1025_inst_req_0;
      type_cast_1025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1025_inst_req_1;
      type_cast_1025_inst_ack_1<= rack(0);
      type_cast_1025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr414_1022,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv417_1026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1035_inst_req_0;
      type_cast_1035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1035_inst_req_1;
      type_cast_1035_inst_ack_1<= rack(0);
      type_cast_1035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr420_1032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv423_1036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_108_inst_req_0;
      type_cast_108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_108_inst_req_1;
      type_cast_108_inst_ack_1<= rack(0);
      type_cast_108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_120_inst_req_0;
      type_cast_120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_120_inst_req_1;
      type_cast_120_inst_ack_1<= rack(0);
      type_cast_120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_133_inst_req_0;
      type_cast_133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_133_inst_req_1;
      type_cast_133_inst_ack_1<= rack(0);
      type_cast_133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_133_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_145_inst_req_0;
      type_cast_145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_145_inst_req_1;
      type_cast_145_inst_ack_1<= rack(0);
      type_cast_145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_158_inst_req_0;
      type_cast_158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_158_inst_req_1;
      type_cast_158_inst_ack_1<= rack(0);
      type_cast_158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1124_155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1125_159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_170_inst_req_0;
      type_cast_170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_170_inst_req_1;
      type_cast_170_inst_ack_1<= rack(0);
      type_cast_170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1128_167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_183_inst_req_0;
      type_cast_183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_183_inst_req_1;
      type_cast_183_inst_ack_1<= rack(0);
      type_cast_183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_193_inst_req_0;
      type_cast_193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_193_inst_req_1;
      type_cast_193_inst_ack_1<= rack(0);
      type_cast_193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inp_d2_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inp_d232_194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_202_inst_req_0;
      type_cast_202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_202_inst_req_1;
      type_cast_202_inst_ack_1<= rack(0);
      type_cast_202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_int_199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_int1_203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inp_d2_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => out_d232_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_220_inst_req_0;
      type_cast_220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_220_inst_req_1;
      type_cast_220_inst_ack_1<= rack(0);
      type_cast_220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out_int_217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => out_int1_221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_265_inst_req_0;
      type_cast_265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_265_inst_req_1;
      type_cast_265_inst_ack_1<= rack(0);
      type_cast_265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp495x_xop_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_288_inst_req_0;
      type_cast_288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_288_inst_req_1;
      type_cast_288_inst_ack_1<= rack(0);
      type_cast_288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext490_439,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_288_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_302_inst_req_0;
      type_cast_302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_302_inst_req_1;
      type_cast_302_inst_ack_1<= rack(0);
      type_cast_302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_315_inst_req_0;
      type_cast_315_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_315_inst_req_1;
      type_cast_315_inst_ack_1<= rack(0);
      type_cast_315_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_316,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_333_inst_req_0;
      type_cast_333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_333_inst_req_1;
      type_cast_333_inst_ack_1<= rack(0);
      type_cast_333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call134_330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_351_inst_req_0;
      type_cast_351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_351_inst_req_1;
      type_cast_351_inst_ack_1<= rack(0);
      type_cast_351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call140_348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv142_352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_369_inst_req_0;
      type_cast_369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_369_inst_req_1;
      type_cast_369_inst_ack_1<= rack(0);
      type_cast_369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_369_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call146_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv148_370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_387_inst_req_0;
      type_cast_387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_387_inst_req_1;
      type_cast_387_inst_ack_1<= rack(0);
      type_cast_387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_405_inst_req_0;
      type_cast_405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_405_inst_req_1;
      type_cast_405_inst_ack_1<= rack(0);
      type_cast_405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call158_402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_423_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_423_inst_req_0;
      type_cast_423_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_423_inst_req_1;
      type_cast_423_inst_ack_1<= rack(0);
      type_cast_423_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_423_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_424,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_45_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_45_inst_req_0;
      type_cast_45_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_45_inst_req_1;
      type_cast_45_inst_ack_1<= rack(0);
      type_cast_45_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_45_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_46,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_485_inst_req_0;
      type_cast_485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_485_inst_req_1;
      type_cast_485_inst_ack_1<= rack(0);
      type_cast_485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp476x_xop_482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_508_inst_req_0;
      type_cast_508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_508_inst_req_1;
      type_cast_508_inst_ack_1<= rack(0);
      type_cast_508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext470_527,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_58_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_58_inst_req_0;
      type_cast_58_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_58_inst_req_1;
      type_cast_58_inst_ack_1<= rack(0);
      type_cast_58_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_58_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_55,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_59,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_631_inst
    process(add_src_597) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_src_597(31 downto 0);
      type_cast_631_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_643_inst
    process(add_out_626) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add_out_626(15 downto 0);
      type_cast_643_wire <= tmp_var; -- 
    end process;
    type_cast_70_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_70_inst_req_0;
      type_cast_70_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_70_inst_req_1;
      type_cast_70_inst_ack_1<= rack(0);
      type_cast_70_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_70_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_71,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_782_inst_req_0;
      type_cast_782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_782_inst_req_1;
      type_cast_782_inst_ack_1<= rack(0);
      type_cast_782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_781_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_787_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_787_inst_req_0;
      type_cast_787_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_787_inst_req_1;
      type_cast_787_inst_ack_1<= rack(0);
      type_cast_787_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_787_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_786_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_797_inst_req_0;
      type_cast_797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_797_inst_req_1;
      type_cast_797_inst_ack_1<= rack(0);
      type_cast_797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_798,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_807_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_807_inst_req_0;
      type_cast_807_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_807_inst_req_1;
      type_cast_807_inst_ack_1<= rack(0);
      type_cast_807_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_807_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr308_804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_808,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr314_814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_827_inst_req_0;
      type_cast_827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_827_inst_req_1;
      type_cast_827_inst_ack_1<= rack(0);
      type_cast_827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_828,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_837_inst_req_0;
      type_cast_837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_837_inst_req_1;
      type_cast_837_inst_ack_1<= rack(0);
      type_cast_837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_80,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_84,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_847_inst_req_1;
      type_cast_847_inst_ack_1<= rack(0);
      type_cast_847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_847_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_857_inst_req_0;
      type_cast_857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_857_inst_req_1;
      type_cast_857_inst_ack_1<= rack(0);
      type_cast_857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_854,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_867_inst_req_0;
      type_cast_867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_867_inst_req_1;
      type_cast_867_inst_ack_1<= rack(0);
      type_cast_867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_867_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_864,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_868,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp464x_xop_924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_111_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_950_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_950_inst_req_0;
      type_cast_950_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_950_inst_req_1;
      type_cast_950_inst_ack_1<= rack(0);
      type_cast_950_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_950_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_950_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_965_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_965_inst_req_0;
      type_cast_965_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_965_inst_req_1;
      type_cast_965_inst_ack_1<= rack(0);
      type_cast_965_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_965_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp377_962,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv381_966,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_975_inst_req_0;
      type_cast_975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_975_inst_req_1;
      type_cast_975_inst_ack_1<= rack(0);
      type_cast_975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr384_972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv387_976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_985_inst_req_0;
      type_cast_985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_985_inst_req_1;
      type_cast_985_inst_ack_1<= rack(0);
      type_cast_985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr390_982,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv393_986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_995_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_995_inst_req_0;
      type_cast_995_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_995_inst_req_1;
      type_cast_995_inst_ack_1<= rack(0);
      type_cast_995_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_995_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr396_992,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv399_996,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_294_index_1_rename
    process(R_indvar489_293_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar489_293_resized;
      ov(13 downto 0) := iv;
      R_indvar489_293_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_294_index_1_resize
    process(indvar489_282) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar489_282;
      ov := iv(13 downto 0);
      R_indvar489_293_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_294_root_address_inst
    process(array_obj_ref_294_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_294_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_294_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_514_index_1_rename
    process(R_indvar469_513_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar469_513_resized;
      ov(13 downto 0) := iv;
      R_indvar469_513_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_514_index_1_resize
    process(indvar469_502) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar469_502;
      ov := iv(13 downto 0);
      R_indvar469_513_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_514_root_address_inst
    process(array_obj_ref_514_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_514_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_514_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_632_index_1_rename
    process(type_cast_631_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_631_resized;
      ov(13 downto 0) := iv;
      type_cast_631_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_632_index_1_resize
    process(type_cast_631_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_631_wire;
      ov := iv(13 downto 0);
      type_cast_631_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_632_root_address_inst
    process(array_obj_ref_632_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_632_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_632_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_644_index_1_rename
    process(type_cast_643_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_643_resized;
      ov(13 downto 0) := iv;
      type_cast_643_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_644_index_1_resize
    process(type_cast_643_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_643_wire;
      ov := iv(13 downto 0);
      type_cast_643_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_644_root_address_inst
    process(array_obj_ref_644_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_644_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_644_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_956_index_1_rename
    process(R_indvar_955_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_955_resized;
      ov(13 downto 0) := iv;
      R_indvar_955_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_956_index_1_resize
    process(indvar_944) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_944;
      ov := iv(13 downto 0);
      R_indvar_955_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_956_root_address_inst
    process(array_obj_ref_956_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_956_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_956_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_addr_0
    process(ptr_deref_431_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_431_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_base_resize
    process(arrayidx_296) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_296;
      ov := iv(13 downto 0);
      ptr_deref_431_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_gather_scatter
    process(add167_429) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add167_429;
      ov(63 downto 0) := iv;
      ptr_deref_431_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_root_address_inst
    process(ptr_deref_431_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_431_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_addr_0
    process(ptr_deref_518_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_518_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_518_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_base_resize
    process(arrayidx269_516) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_516;
      ov := iv(13 downto 0);
      ptr_deref_518_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_gather_scatter
    process(type_cast_520_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_520_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_518_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_root_address_inst
    process(ptr_deref_518_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_518_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_518_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_addr_0
    process(ptr_deref_637_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_637_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_637_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_base_resize
    process(iv1_634) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iv1_634;
      ov := iv(13 downto 0);
      ptr_deref_637_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_gather_scatter
    process(ptr_deref_637_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_637_data_0;
      ov(63 downto 0) := iv;
      i1_638 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_root_address_inst
    process(ptr_deref_637_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_637_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_637_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_651_addr_0
    process(ptr_deref_651_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_651_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_651_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_651_base_resize
    process(ov_647_delayed_6_0_649) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ov_647_delayed_6_0_649;
      ov := iv(13 downto 0);
      ptr_deref_651_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_651_gather_scatter
    process(i1_638) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := i1_638;
      ov(63 downto 0) := iv;
      ptr_deref_651_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_651_root_address_inst
    process(ptr_deref_651_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_651_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_651_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_961_addr_0
    process(ptr_deref_961_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_961_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_961_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_961_base_resize
    process(arrayidx376_958) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx376_958;
      ov := iv(13 downto 0);
      ptr_deref_961_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_961_gather_scatter
    process(ptr_deref_961_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_961_data_0;
      ov(63 downto 0) := iv;
      tmp377_962 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_961_root_address_inst
    process(ptr_deref_961_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_961_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_961_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_575_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_772;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_575_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_575_branch_req_0,
          ack0 => do_while_stmt_575_branch_ack_0,
          ack1 => do_while_stmt_575_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1072_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1071;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1072_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1072_branch_req_0,
          ack0 => if_stmt_1072_branch_ack_0,
          ack1 => if_stmt_1072_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_234_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp467_233;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_234_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_234_branch_req_0,
          ack0 => if_stmt_234_branch_ack_0,
          ack1 => if_stmt_234_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_445_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_444;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_445_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_445_branch_req_0,
          ack0 => if_stmt_445_branch_ack_0,
          ack1 => if_stmt_445_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_458_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264448_457;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_458_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_458_branch_req_0,
          ack0 => if_stmt_458_branch_ack_0,
          ack1 => if_stmt_458_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_533_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_532;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_533_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_533_branch_req_0,
          ack0 => if_stmt_533_branch_ack_0,
          ack1 => if_stmt_533_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_900_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264449_899;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_900_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_900_branch_req_0,
          ack0 => if_stmt_900_branch_ack_0,
          ack1 => if_stmt_900_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_610_inst
    process(nao_606, add_dest_dim1_593) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nao_606, add_dest_dim1_593, tmp_var);
      nao1_611 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_620_inst
    process(input_dim2_585, nao2_616) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_585, nao2_616, tmp_var);
      nao3_621 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_686_inst
    process(input_dim2_585) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_585, konst_685_wire_constant, tmp_var);
      nid2_true_687 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_691_inst
    process(input_dim1_581) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1_581, konst_690_wire_constant, tmp_var);
      nid2_false_692 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_696_inst
    process(add_dest_dim1_593) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim1_593, konst_695_wire_constant, tmp_var);
      nid2_false1_697 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_701_inst
    process(input_dim0_577) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0_577, konst_700_wire_constant, tmp_var);
      nid1_true_702 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_706_inst
    process(add_dest_dim0_589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim0_589, konst_705_wire_constant, tmp_var);
      nid1_true1_707 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_261_inst
    process(tmp495_250) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp495_250, type_cast_260_wire_constant, tmp_var);
      tmp495x_xop_262 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_481_inst
    process(tmp476_470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp476_470, type_cast_480_wire_constant, tmp_var);
      tmp476x_xop_482 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_714_inst
    process(add_src_597) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_src_597, konst_713_wire_constant, tmp_var);
      next_add_src_715 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_923_inst
    process(tmp464_912) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp464_912, type_cast_922_wire_constant, tmp_var);
      tmp464x_xop_924 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1065_inst
    process(indvar_944) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_944, type_cast_1064_wire_constant, tmp_var);
      indvarx_xnext_1066 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_271_inst
    process(iNsTr_19_266) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_19_266, type_cast_270_wire_constant, tmp_var);
      xx_xop503_272 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_438_inst
    process(indvar489_282) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar489_282, type_cast_437_wire_constant, tmp_var);
      indvarx_xnext490_439 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_491_inst
    process(iNsTr_52_486) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_52_486, type_cast_490_wire_constant, tmp_var);
      xx_xop513_492 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_526_inst
    process(indvar469_502) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar469_502, type_cast_525_wire_constant, tmp_var);
      indvarx_xnext470_527 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_933_inst
    process(iNsTr_111_928) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_111_928, type_cast_932_wire_constant, tmp_var);
      xx_xop_934 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_681_inst
    process(NOT_u1_u1_679_wire, cmp_dim1_676) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_679_wire, cmp_dim1_676, tmp_var);
      cmp_dim0_682 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_675_inst
    process(input_dim1_581, SUB_u16_u16_665_665_delayed_1_0_671) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1_581, SUB_u16_u16_665_665_delayed_1_0_671, tmp_var);
      cmp_dim1_676 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1070_inst
    process(indvarx_xnext_1066, tmp468_941) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1066, tmp468_941, tmp_var);
      exitcond1_1071 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_443_inst
    process(indvarx_xnext490_439, tmp500_279) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext490_439, tmp500_279, tmp_var);
      exitcond2_444 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_531_inst
    process(indvarx_xnext470_527, tmp481_499) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext470_527, tmp481_499, tmp_var);
      exitcond_532 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_563_inst
    process(SUB_u16_u16_561_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(SUB_u16_u16_561_wire, konst_562_wire_constant, tmp_var);
      pad_564 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_625_inst
    process(nao3_621) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nao3_621, konst_624_wire_constant, tmp_var);
      add_out_626 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_249_inst
    process(input_size_208) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(input_size_208, type_cast_248_wire_constant, tmp_var);
      tmp495_250 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_469_inst
    process(output_size_226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(output_size_226, type_cast_468_wire_constant, tmp_var);
      tmp476_470 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_911_inst
    process(output_size_226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(output_size_226, type_cast_910_wire_constant, tmp_var);
      tmp464_912 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1001_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_1000_wire_constant, tmp_var);
      shr402_1002 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1011_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_1010_wire_constant, tmp_var);
      shr408_1012 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1021_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_1020_wire_constant, tmp_var);
      shr414_1022 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1031_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_1030_wire_constant, tmp_var);
      shr420_1032 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_803_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_802_wire_constant, tmp_var);
      shr308_804 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_813_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_812_wire_constant, tmp_var);
      shr314_814 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_823_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_822_wire_constant, tmp_var);
      shr320_824 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_833_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_832_wire_constant, tmp_var);
      shr326_834 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_843_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_842_wire_constant, tmp_var);
      shr332_844 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_853_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_852_wire_constant, tmp_var);
      shr338_854 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_863_inst
    process(sub_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_793, type_cast_862_wire_constant, tmp_var);
      shr344_864 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_971_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_970_wire_constant, tmp_var);
      shr384_972 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_981_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_980_wire_constant, tmp_var);
      shr390_982 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_991_inst
    process(tmp377_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_962, type_cast_990_wire_constant, tmp_var);
      shr396_992 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_198_inst
    process(inp_d0_64, inp_d1_89) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(inp_d0_64, inp_d1_89, tmp_var);
      input_int_199 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_216_inst
    process(out_d0_139, out_d1_164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d0_139, out_d1_164, tmp_var);
      out_int_217 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_605_inst
    process(out_d1_164, add_dest_dim0_589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d1_164, add_dest_dim0_589, tmp_var);
      nao_606 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_615_inst
    process(out_d2_189, nao1_611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d2_189, nao1_611, tmp_var);
      nao2_616 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_207_inst
    process(input_int1_203, inp_d232_194) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_int1_203, inp_d232_194, tmp_var);
      input_size_208 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_225_inst
    process(out_int1_221, out_d232_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_int1_221, out_d232_212, tmp_var);
      output_size_226 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_679_inst
    process(cmp_dim2_666) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_666, tmp_var);
      NOT_u1_u1_679_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_721_inst
    process(cmp_dim2_666) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_666, tmp_var);
      NOT_u1_u1_721_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_743_inst
    process(cmp_dim2_666) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_666, tmp_var);
      NOT_u1_u1_743_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_770_inst
    process(cmp_dim0_682) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim0_682, tmp_var);
      NOT_u1_u1_770_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_113_inst
    process(shl18_102, conv20_109) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_102, conv20_109, tmp_var);
      inp_d2_114 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_138_inst
    process(shl114_127, conv116_134) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_127, conv116_134, tmp_var);
      out_d0_139 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_163_inst
    process(shl123_152, conv1125_159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_152, conv1125_159, tmp_var);
      out_d1_164 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_188_inst
    process(shl132_177, conv134_184) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_177, conv134_184, tmp_var);
      out_d2_189 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_63_inst
    process(shl_52, conv3_59) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_52, conv3_59, tmp_var);
      inp_d0_64 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_88_inst
    process(shl9_77, conv11_84) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_77, conv11_84, tmp_var);
      inp_d1_89 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_771_inst
    process(dim0_end_766, NOT_u1_u1_770_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(dim0_end_766, NOT_u1_u1_770_wire, tmp_var);
      continue_flag_772 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_320_inst
    process(shl127_309, conv130_316) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl127_309, conv130_316, tmp_var);
      add131_321 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_338_inst
    process(shl133_327, conv136_334) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl133_327, conv136_334, tmp_var);
      add137_339 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_356_inst
    process(shl139_345, conv142_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl139_345, conv142_352, tmp_var);
      add143_357 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_374_inst
    process(shl145_363, conv148_370) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl145_363, conv148_370, tmp_var);
      add149_375 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_392_inst
    process(shl151_381, conv154_388) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl151_381, conv154_388, tmp_var);
      add155_393 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_410_inst
    process(shl157_399, conv160_406) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl157_399, conv160_406, tmp_var);
      add161_411 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_428_inst
    process(shl163_417, conv166_424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl163_417, conv166_424, tmp_var);
      add167_429 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_101_inst
    process(conv17_96) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_96, type_cast_100_wire_constant, tmp_var);
      shl18_102 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_126_inst
    process(conv113_121) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_121, type_cast_125_wire_constant, tmp_var);
      shl114_127 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_151_inst
    process(conv122_146) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_146, type_cast_150_wire_constant, tmp_var);
      shl123_152 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_176_inst
    process(conv131_171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_171, type_cast_175_wire_constant, tmp_var);
      shl132_177 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_51_inst
    process(conv1_46) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_46, type_cast_50_wire_constant, tmp_var);
      shl_52 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_76_inst
    process(conv8_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_71, type_cast_75_wire_constant, tmp_var);
      shl9_77 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_308_inst
    process(conv125_303) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv125_303, type_cast_307_wire_constant, tmp_var);
      shl127_309 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_326_inst
    process(add131_321) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add131_321, type_cast_325_wire_constant, tmp_var);
      shl133_327 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_344_inst
    process(add137_339) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add137_339, type_cast_343_wire_constant, tmp_var);
      shl139_345 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_362_inst
    process(add143_357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add143_357, type_cast_361_wire_constant, tmp_var);
      shl145_363 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_380_inst
    process(add149_375) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add149_375, type_cast_379_wire_constant, tmp_var);
      shl151_381 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_398_inst
    process(add155_393) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add155_393, type_cast_397_wire_constant, tmp_var);
      shl157_399 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_416_inst
    process(add161_411) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add161_411, type_cast_415_wire_constant, tmp_var);
      shl163_417 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_561_inst
    process(out_d0_139, inp_d0_64) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(out_d0_139, inp_d0_64, tmp_var);
      SUB_u16_u16_561_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_657_inst
    process(inp_d2_114) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(inp_d2_114, konst_656_wire_constant, tmp_var);
      dim2_limit_658 <= tmp_var; --
    end process;
    -- shared split operator group (80) : SUB_u16_u16_670_inst 
    ApIntSub_group_80: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d1_89;
      SUB_u16_u16_665_665_delayed_1_0_671 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_670_inst_req_0;
      SUB_u16_u16_670_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_670_inst_req_1;
      SUB_u16_u16_670_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_80_gI: SplitGuardInterface generic map(name => "ApIntSub_group_80_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_80",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : SUB_u16_u16_760_inst 
    ApIntSub_group_81: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d0_64;
      SUB_u16_u16_749_749_delayed_1_0_761 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_760_inst_req_0;
      SUB_u16_u16_760_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_760_inst_req_1;
      SUB_u16_u16_760_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_81_gI: SplitGuardInterface generic map(name => "ApIntSub_group_81_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_81",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- binary operator SUB_u64_u64_792_inst
    process(conv298_788, conv276_783) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv298_788, conv276_783, tmp_var);
      sub_793 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_231_inst
    process(input_size_208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(input_size_208, type_cast_230_wire_constant, tmp_var);
      cmp467_233 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_255_inst
    process(tmp495_250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp495_250, type_cast_254_wire_constant, tmp_var);
      tmp496_256 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_456_inst
    process(output_size_226) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(output_size_226, type_cast_455_wire_constant, tmp_var);
      cmp264448_457 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_475_inst
    process(tmp476_470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp476_470, type_cast_474_wire_constant, tmp_var);
      tmp477_476 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_898_inst
    process(output_size_226) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(output_size_226, type_cast_897_wire_constant, tmp_var);
      cmp264449_899 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_917_inst
    process(tmp464_912) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp464_912, type_cast_916_wire_constant, tmp_var);
      tmp465_918 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_665_inst
    process(input_dim2_585, dim2_limit_658_delayed_1_0_661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim2_585, dim2_limit_658_delayed_1_0_661, tmp_var);
      cmp_dim2_666 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_765_inst
    process(input_dim0_577, SUB_u16_u16_749_749_delayed_1_0_761) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim0_577, SUB_u16_u16_749_749_delayed_1_0_761, tmp_var);
      dim0_end_766 <= tmp_var; --
    end process;
    -- shared split operator group (91) : array_obj_ref_294_index_offset 
    ApIntAdd_group_91: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar489_293_scaled;
      array_obj_ref_294_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_294_index_offset_req_0;
      array_obj_ref_294_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_294_index_offset_req_1;
      array_obj_ref_294_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_91_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_91_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_91",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : array_obj_ref_514_index_offset 
    ApIntAdd_group_92: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar469_513_scaled;
      array_obj_ref_514_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_514_index_offset_req_0;
      array_obj_ref_514_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_514_index_offset_req_1;
      array_obj_ref_514_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_92_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_92_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_92",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- shared split operator group (93) : array_obj_ref_632_index_offset 
    ApIntAdd_group_93: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_631_scaled;
      array_obj_ref_632_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_632_index_offset_req_0;
      array_obj_ref_632_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_632_index_offset_req_1;
      array_obj_ref_632_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_93_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_93_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_93",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 93
    -- shared split operator group (94) : array_obj_ref_644_index_offset 
    ApIntAdd_group_94: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_643_scaled;
      array_obj_ref_644_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_644_index_offset_req_0;
      array_obj_ref_644_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_644_index_offset_req_1;
      array_obj_ref_644_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_94_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_94_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_94",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 94
    -- shared split operator group (95) : array_obj_ref_956_index_offset 
    ApIntAdd_group_95: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_955_scaled;
      array_obj_ref_956_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_956_index_offset_req_0;
      array_obj_ref_956_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_956_index_offset_req_1;
      array_obj_ref_956_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_95_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_95_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- unary operator type_cast_781_inst
    process(call233_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call233_544, tmp_var);
      type_cast_781_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_786_inst
    process(call297_777) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call297_777, tmp_var);
      type_cast_786_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_637_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_637_load_0_req_0;
      ptr_deref_637_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_637_load_0_req_1;
      ptr_deref_637_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_637_word_address_0;
      ptr_deref_637_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_961_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_961_load_0_req_0;
      ptr_deref_961_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_961_load_0_req_1;
      ptr_deref_961_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_961_word_address_0;
      ptr_deref_961_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_431_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_431_store_0_req_0;
      ptr_deref_431_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_431_store_0_req_1;
      ptr_deref_431_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_431_word_address_0;
      data_in <= ptr_deref_431_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_651_store_0 ptr_deref_518_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_651_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_518_store_0_req_0;
      ptr_deref_651_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_518_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_651_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_518_store_0_req_1;
      ptr_deref_651_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_518_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_651_word_address_0 & ptr_deref_518_word_address_0;
      data_in <= ptr_deref_651_data_0 & ptr_deref_518_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_66_inst RPIPE_ConvTranspose_input_pipe_91_inst RPIPE_ConvTranspose_input_pipe_40_inst RPIPE_ConvTranspose_input_pipe_79_inst RPIPE_ConvTranspose_input_pipe_54_inst RPIPE_ConvTranspose_input_pipe_104_inst RPIPE_ConvTranspose_input_pipe_116_inst RPIPE_ConvTranspose_input_pipe_129_inst RPIPE_ConvTranspose_input_pipe_141_inst RPIPE_ConvTranspose_input_pipe_154_inst RPIPE_ConvTranspose_input_pipe_166_inst RPIPE_ConvTranspose_input_pipe_179_inst RPIPE_ConvTranspose_input_pipe_298_inst RPIPE_ConvTranspose_input_pipe_311_inst RPIPE_ConvTranspose_input_pipe_329_inst RPIPE_ConvTranspose_input_pipe_347_inst RPIPE_ConvTranspose_input_pipe_365_inst RPIPE_ConvTranspose_input_pipe_383_inst RPIPE_ConvTranspose_input_pipe_401_inst RPIPE_ConvTranspose_input_pipe_419_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(159 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 19 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 19 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 19 downto 0);
      signal guard_vector : std_logic_vector( 19 downto 0);
      constant outBUFs : IntegerArray(19 downto 0) := (19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(19 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false);
      constant guardBuffering: IntegerArray(19 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2);
      -- 
    begin -- 
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_79_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_54_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_104_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_129_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_154_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_179_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_311_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_347_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_365_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_383_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_401_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_419_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_79_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_54_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_104_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_129_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_154_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_179_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_311_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_347_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_365_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_383_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_401_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_419_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_79_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_54_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_104_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_129_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_154_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_179_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_311_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_347_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_365_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_383_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_401_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_419_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_79_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_54_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_104_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_129_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_154_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_179_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_311_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_347_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_365_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_383_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_401_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_419_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      call5_67 <= data_out(159 downto 152);
      call14_92 <= data_out(151 downto 144);
      call_41 <= data_out(143 downto 136);
      call10_80 <= data_out(135 downto 128);
      call2_55 <= data_out(127 downto 120);
      call19_105 <= data_out(119 downto 112);
      call110_117 <= data_out(111 downto 104);
      call115_130 <= data_out(103 downto 96);
      call119_142 <= data_out(95 downto 88);
      call1124_155 <= data_out(87 downto 80);
      call1128_167 <= data_out(79 downto 72);
      call133_180 <= data_out(71 downto 64);
      call124_299 <= data_out(63 downto 56);
      call128_312 <= data_out(55 downto 48);
      call134_330 <= data_out(47 downto 40);
      call140_348 <= data_out(39 downto 32);
      call146_366 <= data_out(31 downto 24);
      call152_384 <= data_out(23 downto 16);
      call158_402 <= data_out(15 downto 8);
      call164_420 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 20, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 20,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_872_inst WPIPE_ConvTranspose_output_pipe_869_inst WPIPE_ConvTranspose_output_pipe_878_inst WPIPE_ConvTranspose_output_pipe_875_inst WPIPE_ConvTranspose_output_pipe_884_inst WPIPE_ConvTranspose_output_pipe_881_inst WPIPE_ConvTranspose_output_pipe_1058_inst WPIPE_ConvTranspose_output_pipe_887_inst WPIPE_ConvTranspose_output_pipe_890_inst WPIPE_ConvTranspose_output_pipe_1037_inst WPIPE_ConvTranspose_output_pipe_1049_inst WPIPE_ConvTranspose_output_pipe_1052_inst WPIPE_ConvTranspose_output_pipe_1043_inst WPIPE_ConvTranspose_output_pipe_1046_inst WPIPE_ConvTranspose_output_pipe_1040_inst WPIPE_ConvTranspose_output_pipe_1055_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_872_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_869_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_878_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_875_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_884_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_881_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1058_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_887_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_890_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1037_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1049_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1052_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1043_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1046_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1040_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1055_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_872_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_869_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_878_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_875_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_884_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_881_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1058_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_887_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_890_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1037_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1049_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1052_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1043_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1046_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1040_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1055_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_872_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_869_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_878_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_875_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_884_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_881_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1058_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_887_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_890_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1037_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1049_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1052_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1043_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1046_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1040_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1055_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_872_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_869_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_878_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_875_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_884_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_881_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1058_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_887_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_890_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1037_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1049_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1052_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1043_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1046_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1040_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1055_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv341_858 & conv347_868 & conv329_838 & conv335_848 & conv317_818 & conv323_828 & conv381_966 & conv311_808 & conv305_798 & conv423_1036 & conv399_996 & conv393_986 & conv411_1016 & conv405_1006 & conv417_1026 & conv387_976;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_777_call call_stmt_544_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_777_call_req_0;
      reqL_unguarded(0) <= call_stmt_544_call_req_0;
      call_stmt_777_call_ack_0 <= ackL_unguarded(1);
      call_stmt_544_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_777_call_req_1;
      reqR_unguarded(0) <= call_stmt_544_call_req_1;
      call_stmt_777_call_ack_1 <= ackR_unguarded(1);
      call_stmt_544_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call297_777 <= data_out(127 downto 64);
      call233_544 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad_same_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module zeropad_same
  component zeropad_same is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad_same
  signal zeropad_same_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad_same_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad_same_start_req : std_logic;
  signal zeropad_same_start_ack : std_logic;
  signal zeropad_same_fin_req   : std_logic;
  signal zeropad_same_fin_ack : std_logic;
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(0 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module zeropad_same
  zeropad_same_instance:zeropad_same-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad_same_start_req,
      start_ack => zeropad_same_start_ack,
      fin_req => zeropad_same_fin_req,
      fin_ack => zeropad_same_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad_same_tag_in,
      tag_out => zeropad_same_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad_same_tag_in <= (others => '0');
  zeropad_same_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad_same_start_req, start_ack => zeropad_same_start_ack,  fin_req => zeropad_same_fin_req,  fin_ack => zeropad_same_fin_ack);
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
