-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(63 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_T;
architecture fill_T_arch of fill_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(63 downto 0);
  signal addr_update_enable: Boolean;
  -- output port buffer signals
  signal fill_T_CP_0_start: Boolean;
  signal fill_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_33_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_33_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_37_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_38_inst_req_0 : boolean;
  signal CONCAT_u8_u16_38_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_38_inst_req_1 : boolean;
  signal CONCAT_u8_u16_38_inst_ack_1 : boolean;
  signal CONCAT_u48_u64_45_inst_req_0 : boolean;
  signal CONCAT_u48_u64_45_inst_ack_0 : boolean;
  signal CONCAT_u48_u64_45_inst_req_1 : boolean;
  signal CONCAT_u48_u64_45_inst_ack_1 : boolean;
  signal if_stmt_47_branch_req_0 : boolean;
  signal if_stmt_47_branch_ack_1 : boolean;
  signal if_stmt_47_branch_ack_0 : boolean;
  signal phi_stmt_15_req_1 : boolean;
  signal phi_stmt_21_req_0 : boolean;
  signal nmycount_31_17_buf_req_0 : boolean;
  signal nmycount_31_17_buf_ack_0 : boolean;
  signal nmycount_31_17_buf_req_1 : boolean;
  signal nmycount_31_17_buf_ack_1 : boolean;
  signal phi_stmt_15_req_0 : boolean;
  signal ninput_word_46_25_buf_req_0 : boolean;
  signal ninput_word_46_25_buf_ack_0 : boolean;
  signal ninput_word_46_25_buf_req_1 : boolean;
  signal ninput_word_46_25_buf_ack_1 : boolean;
  signal phi_stmt_21_req_1 : boolean;
  signal phi_stmt_15_ack_0 : boolean;
  signal phi_stmt_21_ack_0 : boolean;
  signal array_obj_ref_60_index_offset_req_0 : boolean;
  signal array_obj_ref_60_index_offset_ack_0 : boolean;
  signal array_obj_ref_60_index_offset_req_1 : boolean;
  signal array_obj_ref_60_index_offset_ack_1 : boolean;
  signal addr_of_61_final_reg_req_0 : boolean;
  signal addr_of_61_final_reg_ack_0 : boolean;
  signal addr_of_61_final_reg_req_1 : boolean;
  signal addr_of_61_final_reg_ack_1 : boolean;
  signal ptr_deref_64_store_0_req_0 : boolean;
  signal ptr_deref_64_store_0_ack_0 : boolean;
  signal ptr_deref_64_store_0_req_1 : boolean;
  signal ptr_deref_64_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_T_CP_0: Block -- control-path 
    signal fill_T_CP_0_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    fill_T_CP_0_elements(0) <= fill_T_CP_0_start;
    fill_T_CP_0_symbol <= fill_T_CP_0_elements(33);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_13/$entry
      -- CP-element group 0: 	 branch_block_stmt_13/branch_block_stmt_13__entry__
      -- CP-element group 0: 	 branch_block_stmt_13/merge_stmt_14__entry__
      -- CP-element group 0: 	 branch_block_stmt_13/merge_stmt_14_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	26 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	2 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (12) 
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_update_start_
      -- CP-element group 1: 	 branch_block_stmt_13/merge_stmt_14__exit__
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46__entry__
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_update_start_
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Update/cr
      -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => RPIPE_maxpool_input_pipe_33_inst_req_0); -- 
    cr_57_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_57_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u8_u16_38_inst_req_1); -- 
    cr_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u48_u64_45_inst_req_1); -- 
    fill_T_CP_0_elements(1) <= fill_T_CP_0_elements(26);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_update_start_
      -- CP-element group 2: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Sample/$exit
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_33_inst_ack_0, ack => fill_T_CP_0_elements(2)); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(2), ack => RPIPE_maxpool_input_pipe_33_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_33_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/rr
      -- 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_33_inst_ack_1, ack => fill_T_CP_0_elements(3)); -- 
    rr_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(3), ack => RPIPE_maxpool_input_pipe_37_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_update_start_
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/cr
      -- 
    ra_43_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_37_inst_ack_0, ack => fill_T_CP_0_elements(4)); -- 
    cr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(4), ack => RPIPE_maxpool_input_pipe_37_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/RPIPE_maxpool_input_pipe_37_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/rr
      -- 
    ca_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_37_inst_ack_1, ack => fill_T_CP_0_elements(5)); -- 
    rr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(5), ack => CONCAT_u8_u16_38_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Sample/ra
      -- 
    ra_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_38_inst_ack_0, ack => fill_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u8_u16_38_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Sample/rr
      -- 
    ca_58_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_38_inst_ack_1, ack => fill_T_CP_0_elements(7)); -- 
    rr_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => CONCAT_u48_u64_45_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Sample/ra
      -- 
    ra_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u48_u64_45_inst_ack_0, ack => fill_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (27) 
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46__exit__
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47__entry__
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/assign_stmt_31_to_assign_stmt_46/CONCAT_u48_u64_45_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/ULT_u4_u1_50_inputs/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/ULT_u4_u1_50_inputs/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/cr
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/ULT_u4_u1_50/SplitProtocol/Update/ca
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_13/ULT_u4_u1_50_place
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_13/if_stmt_47_else_link/$entry
      -- 
    ca_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u48_u64_45_inst_ack_1, ack => fill_T_CP_0_elements(9)); -- 
    branch_req_99_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_99_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(9), ack => if_stmt_47_branch_req_0); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	20 
    -- CP-element group 10:  members (18) 
      -- CP-element group 10: 	 branch_block_stmt_13/if_stmt_47_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_13/if_stmt_47_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_13/loopback
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/req
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/req
      -- 
    if_choice_transition_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_47_branch_ack_1, ack => fill_T_CP_0_elements(10)); -- 
    req_148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => nmycount_31_17_buf_req_0); -- 
    req_153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => nmycount_31_17_buf_req_1); -- 
    req_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => ninput_word_46_25_buf_req_0); -- 
    req_173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => ninput_word_46_25_buf_req_1); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	27 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	30 
    -- CP-element group 11: 	32 
    -- CP-element group 11:  members (30) 
      -- CP-element group 11: 	 branch_block_stmt_13/$exit
      -- CP-element group 11: 	 branch_block_stmt_13/branch_block_stmt_13__exit__
      -- CP-element group 11: 	 branch_block_stmt_13/if_stmt_47__exit__
      -- CP-element group 11: 	 branch_block_stmt_13/if_stmt_47_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_13/if_stmt_47_else_link/else_choice_transition
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_update_start_
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resized_1
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scaled_1
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_computed_1
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/$exit
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/index_resize_req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_resize_1/index_resize_ack
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/$exit
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/scale_rename_req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_index_scale_1/scale_rename_ack
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_update_start
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/req
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_update_start_
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_47_branch_ack_0, ack => fill_T_CP_0_elements(11)); -- 
    req_209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => array_obj_ref_60_index_offset_req_0); -- 
    req_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => array_obj_ref_60_index_offset_req_1); -- 
    req_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => addr_of_61_final_reg_req_1); -- 
    cr_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => ptr_deref_64_store_0_req_1); -- 
    -- CP-element group 12:  fork  transition  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_sources/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/$entry
      -- CP-element group 12: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_sources/$entry
      -- 
    fill_T_CP_0_elements(12) <= fill_T_CP_0_elements(0);
    -- CP-element group 13:  transition  output  delay-element  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/$exit
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_sources/$exit
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_sources/type_cast_20_konst_delay_trans
      -- CP-element group 13: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_15/phi_stmt_15_req
      -- 
    phi_stmt_15_req_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15_req_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(13), ack => phi_stmt_15_req_1); -- 
    -- Element group fill_T_CP_0_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(12), ack => fill_T_CP_0_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  transition  output  delay-element  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/$exit
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_sources/type_cast_24_konst_delay_trans
      -- CP-element group 14: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/phi_stmt_21/phi_stmt_21_req
      -- 
    phi_stmt_21_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_21_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => phi_stmt_21_req_0); -- 
    -- Element group fill_T_CP_0_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(12), ack => fill_T_CP_0_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  transition  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	23 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_13/merge_stmt_14__entry___PhiReq/$exit
      -- 
    fill_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(13) & fill_T_CP_0_elements(14);
      gj_fill_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Sample/ack
      -- 
    ack_149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_31_17_buf_ack_0, ack => fill_T_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/Update/ack
      -- 
    ack_154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_31_17_buf_ack_1, ack => fill_T_CP_0_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/$exit
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/$exit
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_sources/Interlock/$exit
      -- CP-element group 18: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_15/phi_stmt_15_req
      -- 
    phi_stmt_15_req_155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15_req_155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(18), ack => phi_stmt_15_req_0); -- 
    fill_T_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(16) & fill_T_CP_0_elements(17);
      gj_fill_T_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Sample/ack
      -- 
    ack_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_46_25_buf_ack_0, ack => fill_T_CP_0_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/Update/ack
      -- 
    ack_174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_46_25_buf_ack_1, ack => fill_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/$exit
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/$exit
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_sources/Interlock/$exit
      -- CP-element group 21: 	 branch_block_stmt_13/loopback_PhiReq/phi_stmt_21/phi_stmt_21_req
      -- 
    phi_stmt_21_req_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_21_req_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(21), ack => phi_stmt_21_req_1); -- 
    fill_T_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(19) & fill_T_CP_0_elements(20);
      gj_fill_T_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_13/loopback_PhiReq/$exit
      -- 
    fill_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(18) & fill_T_CP_0_elements(21);
      gj_fill_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  merge  fork  transition  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_13/merge_stmt_14_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/$entry
      -- 
    fill_T_CP_0_elements(23) <= OrReduce(fill_T_CP_0_elements(15) & fill_T_CP_0_elements(22));
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/phi_stmt_15_ack
      -- 
    phi_stmt_15_ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_15_ack_0, ack => fill_T_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/phi_stmt_21_ack
      -- 
    phi_stmt_21_ack_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_21_ack_0, ack => fill_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	1 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_13/merge_stmt_14_PhiAck/$exit
      -- 
    fill_T_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(24) & fill_T_CP_0_elements(25);
      gj_fill_T_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	11 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_sample_complete
      -- CP-element group 27: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Sample/ack
      -- 
    ack_210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_60_index_offset_ack_0, ack => fill_T_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	11 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (11) 
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_sample_start_
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_offset_calculated
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/$exit
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/array_obj_ref_60_final_index_sum_regn_Update/ack
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/$entry
      -- CP-element group 28: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/req
      -- 
    ack_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_60_index_offset_ack_1, ack => fill_T_CP_0_elements(28)); -- 
    req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(28), ack => addr_of_61_final_reg_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_sample_completed_
      -- CP-element group 29: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/$exit
      -- CP-element group 29: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_request/ack
      -- 
    ack_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_61_final_reg_ack_0, ack => fill_T_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	11 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (28) 
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_update_completed_
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/addr_of_61_complete/ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_sample_start_
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_address_calculated
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_address_calculated
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_root_address_calculated
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_address_resized
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/base_resize_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_addr_resize/base_resize_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/root_register_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_word_addrgen/root_register_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/$exit
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/split_req
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/ptr_deref_64_Split/split_ack
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/rr
      -- 
    ack_230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_61_final_reg_ack_1, ack => fill_T_CP_0_elements(30)); -- 
    rr_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(30), ack => ptr_deref_64_store_0_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_sample_completed_
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/$exit
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Sample/word_access_start/word_0/ra
      -- 
    ra_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_64_store_0_ack_0, ack => fill_T_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	11 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_update_completed_
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/$exit
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/$exit
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_62_to_assign_stmt_66/ptr_deref_64_Update/word_access_complete/word_0/ca
      -- 
    ca_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_64_store_0_ack_1, ack => fill_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 $exit
      -- CP-element group 33: 	 assign_stmt_62_to_assign_stmt_66/$exit
      -- 
    fill_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(27) & fill_T_CP_0_elements(32);
      gj_fill_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_maxpool_input_pipe_37_wire : std_logic_vector(7 downto 0);
    signal R_addr_59_resized : std_logic_vector(13 downto 0);
    signal R_addr_59_scaled : std_logic_vector(13 downto 0);
    signal ULT_u4_u1_50_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_60_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_60_root_address : std_logic_vector(13 downto 0);
    signal input_word_21 : std_logic_vector(63 downto 0);
    signal konst_29_wire_constant : std_logic_vector(3 downto 0);
    signal konst_49_wire_constant : std_logic_vector(3 downto 0);
    signal mycount_15 : std_logic_vector(3 downto 0);
    signal ninput_word_46 : std_logic_vector(63 downto 0);
    signal ninput_word_46_25_buffered : std_logic_vector(63 downto 0);
    signal nmycount_31 : std_logic_vector(3 downto 0);
    signal nmycount_31_17_buffered : std_logic_vector(3 downto 0);
    signal ptr_62 : std_logic_vector(31 downto 0);
    signal ptr_deref_64_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_64_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_64_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_64_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_64_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_64_word_offset_0 : std_logic_vector(13 downto 0);
    signal slice_43_wire : std_logic_vector(47 downto 0);
    signal type_cast_20_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_24_wire_constant : std_logic_vector(63 downto 0);
    signal val1_34 : std_logic_vector(7 downto 0);
    signal val_39 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_60_constant_part_of_offset <= "00000000000000";
    array_obj_ref_60_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_60_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_60_resized_base_address <= "00000000000000";
    konst_29_wire_constant <= "0001";
    konst_49_wire_constant <= "0011";
    ptr_deref_64_word_offset_0 <= "00000000000000";
    type_cast_20_wire_constant <= "0000";
    type_cast_24_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_15: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_31_17_buffered & type_cast_20_wire_constant;
      req <= phi_stmt_15_req_0 & phi_stmt_15_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_15",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_15_ack_0,
          idata => idata,
          odata => mycount_15,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_15
    phi_stmt_21: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_24_wire_constant & ninput_word_46_25_buffered;
      req <= phi_stmt_21_req_0 & phi_stmt_21_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_21",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_21_ack_0,
          idata => idata,
          odata => input_word_21,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_21
    -- flow-through slice operator slice_43_inst
    slice_43_wire <= input_word_21(47 downto 0);
    addr_of_61_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_61_final_reg_req_0;
      addr_of_61_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_61_final_reg_req_1;
      addr_of_61_final_reg_ack_1<= rack(0);
      addr_of_61_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_61_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_60_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_62,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ninput_word_46_25_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ninput_word_46_25_buf_req_0;
      ninput_word_46_25_buf_ack_0<= wack(0);
      rreq(0) <= ninput_word_46_25_buf_req_1;
      ninput_word_46_25_buf_ack_1<= rack(0);
      ninput_word_46_25_buf : InterlockBuffer generic map ( -- 
        name => "ninput_word_46_25_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ninput_word_46,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ninput_word_46_25_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_31_17_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_31_17_buf_req_0;
      nmycount_31_17_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_31_17_buf_req_1;
      nmycount_31_17_buf_ack_1<= rack(0);
      nmycount_31_17_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_31_17_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_31,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_31_17_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_60_index_1_rename
    process(R_addr_59_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_59_resized;
      ov(13 downto 0) := iv;
      R_addr_59_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_59_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_60_root_address_inst
    process(array_obj_ref_60_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_60_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_60_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_addr_0
    process(ptr_deref_64_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_64_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_64_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_base_resize
    process(ptr_62) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_62;
      ov := iv(13 downto 0);
      ptr_deref_64_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_gather_scatter
    process(ninput_word_46) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ninput_word_46;
      ov(63 downto 0) := iv;
      ptr_deref_64_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_64_root_address_inst
    process(ptr_deref_64_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_64_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_64_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_47_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u4_u1_50_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_47_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_47_branch_req_0,
          ack0 => if_stmt_47_branch_ack_0,
          ack1 => if_stmt_47_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u4_u4_30_inst
    process(mycount_15) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_15, konst_29_wire_constant, tmp_var);
      nmycount_31 <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u48_u64_45_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_43_wire & val_39;
      ninput_word_46 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u48_u64_45_inst_req_0;
      CONCAT_u48_u64_45_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u48_u64_45_inst_req_1;
      CONCAT_u48_u64_45_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 48,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : CONCAT_u8_u16_38_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= val1_34 & RPIPE_maxpool_input_pipe_37_wire;
      val_39 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u8_u16_38_inst_req_0;
      CONCAT_u8_u16_38_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_38_inst_req_1;
      CONCAT_u8_u16_38_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator ULT_u4_u1_50_inst
    process(mycount_15) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_15, konst_49_wire_constant, tmp_var);
      ULT_u4_u1_50_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : array_obj_ref_60_index_offset 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_59_scaled;
      array_obj_ref_60_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_60_index_offset_req_0;
      array_obj_ref_60_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_60_index_offset_req_1;
      array_obj_ref_60_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared store operator group (0) : ptr_deref_64_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_64_store_0_req_0;
      ptr_deref_64_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_64_store_0_req_1;
      ptr_deref_64_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_64_word_address_0;
      data_in <= ptr_deref_64_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_33_inst RPIPE_maxpool_input_pipe_37_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_33_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_37_inst_req_0;
      RPIPE_maxpool_input_pipe_33_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_37_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_33_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_37_inst_req_1;
      RPIPE_maxpool_input_pipe_33_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_37_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      val1_34 <= data_out(15 downto 8);
      RPIPE_maxpool_input_pipe_37_wire <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end fill_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    fill_T_call_reqs : out  std_logic_vector(0 downto 0);
    fill_T_call_acks : in   std_logic_vector(0 downto 0);
    fill_T_call_data : out  std_logic_vector(63 downto 0);
    fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_T_return_reqs : out  std_logic_vector(0 downto 0);
    fill_T_return_acks : in   std_logic_vector(0 downto 0);
    fill_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_call_acks : in   std_logic_vector(0 downto 0);
    maxPool4_call_data : out  std_logic_vector(159 downto 0);
    maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
    maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_return_acks : in   std_logic_vector(0 downto 0);
    maxPool4_return_data : in   std_logic_vector(7 downto 0);
    maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(31 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool3D;
architecture maxPool3D_arch of maxPool3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal maxPool3D_CP_1610_start: Boolean;
  signal maxPool3D_CP_1610_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_685_inst_req_0 : boolean;
  signal type_cast_652_inst_ack_0 : boolean;
  signal type_cast_639_inst_ack_1 : boolean;
  signal type_cast_677_inst_req_0 : boolean;
  signal type_cast_906_inst_ack_0 : boolean;
  signal type_cast_652_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_610_inst_ack_1 : boolean;
  signal type_cast_589_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_660_inst_req_0 : boolean;
  signal type_cast_627_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_610_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_623_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_685_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_req_0 : boolean;
  signal type_cast_639_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_610_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_635_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_660_inst_ack_1 : boolean;
  signal type_cast_589_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_610_inst_req_1 : boolean;
  signal type_cast_589_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_ack_0 : boolean;
  signal type_cast_664_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_635_inst_req_1 : boolean;
  signal type_cast_589_inst_ack_0 : boolean;
  signal type_cast_639_inst_req_1 : boolean;
  signal type_cast_627_inst_ack_1 : boolean;
  signal type_cast_652_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_660_inst_ack_0 : boolean;
  signal type_cast_639_inst_req_0 : boolean;
  signal type_cast_677_inst_ack_1 : boolean;
  signal type_cast_1025_inst_req_0 : boolean;
  signal type_cast_906_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_673_inst_req_0 : boolean;
  signal type_cast_911_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_673_inst_ack_0 : boolean;
  signal type_cast_911_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_673_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_673_inst_ack_1 : boolean;
  signal type_cast_602_inst_req_0 : boolean;
  signal call_stmt_987_call_ack_0 : boolean;
  signal call_stmt_987_call_req_0 : boolean;
  signal type_cast_602_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_req_1 : boolean;
  signal type_cast_677_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_685_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_635_inst_req_0 : boolean;
  signal type_cast_664_inst_req_0 : boolean;
  signal type_cast_652_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_585_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_660_inst_req_1 : boolean;
  signal type_cast_664_inst_req_1 : boolean;
  signal type_cast_614_inst_req_0 : boolean;
  signal type_cast_614_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_585_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_635_inst_ack_0 : boolean;
  signal type_cast_602_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_598_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_585_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_585_inst_ack_0 : boolean;
  signal type_cast_602_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_598_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_623_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_623_inst_req_0 : boolean;
  signal type_cast_614_inst_req_1 : boolean;
  signal type_cast_627_inst_req_0 : boolean;
  signal type_cast_614_inst_ack_1 : boolean;
  signal type_cast_627_inst_ack_0 : boolean;
  signal type_cast_677_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_623_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_685_inst_ack_1 : boolean;
  signal type_cast_664_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_598_inst_req_1 : boolean;
  signal call_stmt_987_call_req_1 : boolean;
  signal call_stmt_987_call_ack_1 : boolean;
  signal type_cast_906_inst_ack_1 : boolean;
  signal type_cast_911_inst_req_1 : boolean;
  signal type_cast_1083_inst_req_0 : boolean;
  signal type_cast_911_inst_ack_1 : boolean;
  signal call_stmt_1100_call_req_1 : boolean;
  signal if_stmt_1053_branch_ack_1 : boolean;
  signal call_stmt_1066_call_req_0 : boolean;
  signal type_cast_1083_inst_ack_0 : boolean;
  signal call_stmt_1100_call_ack_1 : boolean;
  signal call_stmt_1066_call_ack_0 : boolean;
  signal call_stmt_1066_call_req_1 : boolean;
  signal if_stmt_1053_branch_ack_0 : boolean;
  signal type_cast_1001_inst_req_0 : boolean;
  signal type_cast_1001_inst_ack_0 : boolean;
  signal type_cast_1025_inst_ack_0 : boolean;
  signal type_cast_1001_inst_req_1 : boolean;
  signal type_cast_1001_inst_ack_1 : boolean;
  signal type_cast_1083_inst_req_1 : boolean;
  signal call_stmt_1066_call_ack_1 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1077_inst_req_0 : boolean;
  signal W_colx_x1_1002_delayed_1_0_1003_inst_req_0 : boolean;
  signal W_colx_x1_1002_delayed_1_0_1003_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1077_inst_ack_0 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal type_cast_1025_inst_req_1 : boolean;
  signal W_colx_x1_1002_delayed_1_0_1003_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_598_inst_ack_1 : boolean;
  signal type_cast_689_inst_req_0 : boolean;
  signal if_stmt_1053_branch_req_0 : boolean;
  signal type_cast_689_inst_ack_0 : boolean;
  signal type_cast_689_inst_req_1 : boolean;
  signal type_cast_689_inst_ack_1 : boolean;
  signal type_cast_1070_inst_ack_1 : boolean;
  signal type_cast_1070_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_698_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_698_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_698_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_698_inst_ack_1 : boolean;
  signal call_stmt_1100_call_ack_0 : boolean;
  signal type_cast_924_inst_ack_1 : boolean;
  signal type_cast_924_inst_req_1 : boolean;
  signal type_cast_702_inst_req_0 : boolean;
  signal type_cast_702_inst_ack_0 : boolean;
  signal type_cast_1087_inst_ack_1 : boolean;
  signal type_cast_702_inst_req_1 : boolean;
  signal type_cast_702_inst_ack_1 : boolean;
  signal type_cast_1070_inst_ack_0 : boolean;
  signal type_cast_1070_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_710_inst_req_0 : boolean;
  signal do_while_stmt_896_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_710_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_710_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_710_inst_ack_1 : boolean;
  signal call_stmt_1100_call_req_0 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal type_cast_714_inst_req_0 : boolean;
  signal do_while_stmt_896_branch_ack_0 : boolean;
  signal type_cast_714_inst_ack_0 : boolean;
  signal type_cast_1087_inst_req_1 : boolean;
  signal type_cast_714_inst_req_1 : boolean;
  signal type_cast_714_inst_ack_1 : boolean;
  signal type_cast_1062_inst_ack_1 : boolean;
  signal type_cast_1062_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_723_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_723_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_723_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_723_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal W_rowx_x1_1023_delayed_2_0_1027_inst_ack_1 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal W_rowx_x1_1023_delayed_2_0_1027_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal phi_stmt_908_ack_0 : boolean;
  signal type_cast_906_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1077_inst_ack_1 : boolean;
  signal type_cast_920_inst_ack_1 : boolean;
  signal type_cast_920_inst_req_1 : boolean;
  signal type_cast_737_inst_req_0 : boolean;
  signal type_cast_737_inst_ack_0 : boolean;
  signal type_cast_1087_inst_ack_0 : boolean;
  signal type_cast_737_inst_req_1 : boolean;
  signal W_rowx_x1_1023_delayed_2_0_1027_inst_ack_0 : boolean;
  signal type_cast_737_inst_ack_1 : boolean;
  signal type_cast_1062_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1077_inst_req_1 : boolean;
  signal type_cast_1087_inst_req_0 : boolean;
  signal phi_stmt_908_req_1 : boolean;
  signal if_stmt_755_branch_req_0 : boolean;
  signal type_cast_920_inst_ack_0 : boolean;
  signal if_stmt_755_branch_ack_1 : boolean;
  signal if_stmt_755_branch_ack_0 : boolean;
  signal W_rowx_x1_1023_delayed_2_0_1027_inst_req_0 : boolean;
  signal type_cast_920_inst_req_0 : boolean;
  signal type_cast_792_inst_req_0 : boolean;
  signal type_cast_792_inst_ack_0 : boolean;
  signal type_cast_792_inst_req_1 : boolean;
  signal type_cast_792_inst_ack_1 : boolean;
  signal type_cast_1062_inst_req_0 : boolean;
  signal call_stmt_818_call_req_0 : boolean;
  signal call_stmt_818_call_ack_0 : boolean;
  signal call_stmt_818_call_req_1 : boolean;
  signal call_stmt_818_call_ack_1 : boolean;
  signal phi_stmt_908_req_0 : boolean;
  signal if_stmt_830_branch_req_0 : boolean;
  signal W_colx_x1_1002_delayed_1_0_1003_inst_ack_1 : boolean;
  signal if_stmt_830_branch_ack_1 : boolean;
  signal if_stmt_830_branch_ack_0 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal call_stmt_853_call_req_0 : boolean;
  signal type_cast_1025_inst_ack_1 : boolean;
  signal call_stmt_853_call_ack_0 : boolean;
  signal call_stmt_853_call_req_1 : boolean;
  signal call_stmt_853_call_ack_1 : boolean;
  signal type_cast_857_inst_req_0 : boolean;
  signal type_cast_857_inst_ack_0 : boolean;
  signal type_cast_857_inst_req_1 : boolean;
  signal type_cast_857_inst_ack_1 : boolean;
  signal type_cast_861_inst_req_0 : boolean;
  signal type_cast_861_inst_ack_0 : boolean;
  signal type_cast_861_inst_req_1 : boolean;
  signal type_cast_861_inst_ack_1 : boolean;
  signal type_cast_865_inst_req_0 : boolean;
  signal type_cast_865_inst_ack_0 : boolean;
  signal type_cast_865_inst_req_1 : boolean;
  signal type_cast_865_inst_ack_1 : boolean;
  signal do_while_stmt_896_branch_req_0 : boolean;
  signal phi_stmt_898_req_0 : boolean;
  signal phi_stmt_898_req_1 : boolean;
  signal phi_stmt_898_ack_0 : boolean;
  signal type_cast_1083_inst_ack_1 : boolean;
  signal type_cast_901_inst_req_0 : boolean;
  signal type_cast_901_inst_ack_0 : boolean;
  signal type_cast_901_inst_req_1 : boolean;
  signal type_cast_901_inst_ack_1 : boolean;
  signal phi_stmt_903_req_0 : boolean;
  signal phi_stmt_903_req_1 : boolean;
  signal phi_stmt_903_ack_0 : boolean;
  signal phi_stmt_809_req_0 : boolean;
  signal type_cast_815_inst_req_0 : boolean;
  signal type_cast_815_inst_ack_0 : boolean;
  signal type_cast_815_inst_req_1 : boolean;
  signal type_cast_815_inst_ack_1 : boolean;
  signal phi_stmt_809_req_1 : boolean;
  signal phi_stmt_809_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool3D_CP_1610_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_1610_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool3D_CP_1610_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_1610_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool3D_CP_1610: Block -- control-path 
    signal maxPool3D_CP_1610_elements: BooleanArray(204 downto 0);
    -- 
  begin -- 
    maxPool3D_CP_1610_elements(0) <= maxPool3D_CP_1610_start;
    maxPool3D_CP_1610_symbol <= maxPool3D_CP_1610_elements(197);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (44) 
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_583/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/branch_block_stmt_583__entry__
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733__entry__
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_update_start_
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Update/cr
      -- 
    cr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_589_inst_req_1); -- 
    cr_1773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_627_inst_req_1); -- 
    cr_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_639_inst_req_1); -- 
    cr_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_652_inst_req_1); -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => RPIPE_maxpool_input_pipe_585_inst_req_0); -- 
    cr_1857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_664_inst_req_1); -- 
    cr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_602_inst_req_1); -- 
    cr_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_614_inst_req_1); -- 
    cr_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_677_inst_req_1); -- 
    cr_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_689_inst_req_1); -- 
    cr_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_702_inst_req_1); -- 
    cr_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_714_inst_req_1); -- 
    cr_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(0), ack => type_cast_727_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	180 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	181 
    -- CP-element group 1: 	182 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_583/do_while_stmt_896__exit__
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053__entry__
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_583/if_stmt_1053_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_583/R_whilex_xbody_whilex_xend_taken_1054_place
      -- 
    branch_req_2434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(1), ack => if_stmt_1053_branch_req_0); -- 
    maxPool3D_CP_1610_elements(1) <= maxPool3D_CP_1610_elements(180);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_update_start_
      -- CP-element group 2: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Update/$entry
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_585_inst_ack_0, ack => maxPool3D_CP_1610_elements(2)); -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(2), ack => RPIPE_maxpool_input_pipe_585_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_585_Update/ca
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_585_inst_ack_1, ack => maxPool3D_CP_1610_elements(3)); -- 
    rr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(3), ack => type_cast_589_inst_req_0); -- 
    rr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(3), ack => RPIPE_maxpool_input_pipe_598_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Sample/$exit
      -- 
    ra_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_589_inst_ack_0, ack => maxPool3D_CP_1610_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_589_Update/ca
      -- 
    ca_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_589_inst_ack_1, ack => maxPool3D_CP_1610_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_update_start_
      -- CP-element group 6: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Update/cr
      -- 
    ra_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_598_inst_ack_0, ack => maxPool3D_CP_1610_elements(6)); -- 
    cr_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(6), ack => RPIPE_maxpool_input_pipe_598_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_598_Update/ca
      -- 
    ca_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_598_inst_ack_1, ack => maxPool3D_CP_1610_elements(7)); -- 
    rr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(7), ack => type_cast_602_inst_req_0); -- 
    rr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(7), ack => RPIPE_maxpool_input_pipe_610_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Sample/ra
      -- 
    ra_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_602_inst_ack_0, ack => maxPool3D_CP_1610_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_602_Update/ca
      -- 
    ca_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_602_inst_ack_1, ack => maxPool3D_CP_1610_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_update_start_
      -- CP-element group 10: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_sample_completed_
      -- 
    ra_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_610_inst_ack_0, ack => maxPool3D_CP_1610_elements(10)); -- 
    cr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(10), ack => RPIPE_maxpool_input_pipe_610_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_610_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_sample_start_
      -- 
    ca_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_610_inst_ack_1, ack => maxPool3D_CP_1610_elements(11)); -- 
    rr_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(11), ack => type_cast_614_inst_req_0); -- 
    rr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(11), ack => RPIPE_maxpool_input_pipe_623_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Sample/ra
      -- 
    ra_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_0, ack => maxPool3D_CP_1610_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	50 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_614_Update/ca
      -- 
    ca_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_1, ack => maxPool3D_CP_1610_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_update_start_
      -- CP-element group 14: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Sample/ra
      -- 
    ra_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_623_inst_ack_0, ack => maxPool3D_CP_1610_elements(14)); -- 
    cr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(14), ack => RPIPE_maxpool_input_pipe_623_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_623_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_sample_start_
      -- 
    ca_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_623_inst_ack_1, ack => maxPool3D_CP_1610_elements(15)); -- 
    rr_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(15), ack => type_cast_627_inst_req_0); -- 
    rr_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(15), ack => RPIPE_maxpool_input_pipe_635_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Sample/ra
      -- 
    ra_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_0, ack => maxPool3D_CP_1610_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	50 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_627_Update/ca
      -- 
    ca_1774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_1, ack => maxPool3D_CP_1610_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_update_start_
      -- CP-element group 18: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Sample/ra
      -- 
    ra_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_635_inst_ack_0, ack => maxPool3D_CP_1610_elements(18)); -- 
    cr_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(18), ack => RPIPE_maxpool_input_pipe_635_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_635_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Sample/$entry
      -- 
    ca_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_635_inst_ack_1, ack => maxPool3D_CP_1610_elements(19)); -- 
    rr_1796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(19), ack => type_cast_639_inst_req_0); -- 
    rr_1810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(19), ack => RPIPE_maxpool_input_pipe_648_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Sample/$exit
      -- 
    ra_1797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_0, ack => maxPool3D_CP_1610_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	50 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_639_Update/$exit
      -- 
    ca_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_1, ack => maxPool3D_CP_1610_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_update_start_
      -- CP-element group 22: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Sample/$exit
      -- 
    ra_1811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_648_inst_ack_0, ack => maxPool3D_CP_1610_elements(22)); -- 
    cr_1815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(22), ack => RPIPE_maxpool_input_pipe_648_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_648_Update/ca
      -- 
    ca_1816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_648_inst_ack_1, ack => maxPool3D_CP_1610_elements(23)); -- 
    rr_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(23), ack => RPIPE_maxpool_input_pipe_660_inst_req_0); -- 
    rr_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(23), ack => type_cast_652_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_sample_completed_
      -- 
    ra_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_0, ack => maxPool3D_CP_1610_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_652_Update/ca
      -- 
    ca_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_1, ack => maxPool3D_CP_1610_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_update_start_
      -- 
    ra_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_660_inst_ack_0, ack => maxPool3D_CP_1610_elements(26)); -- 
    cr_1843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(26), ack => RPIPE_maxpool_input_pipe_660_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_660_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_sample_start_
      -- 
    ca_1844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_660_inst_ack_1, ack => maxPool3D_CP_1610_elements(27)); -- 
    rr_1852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(27), ack => type_cast_664_inst_req_0); -- 
    rr_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(27), ack => RPIPE_maxpool_input_pipe_673_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Sample/$exit
      -- 
    ra_1853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_0, ack => maxPool3D_CP_1610_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	50 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_664_Update/ca
      -- 
    ca_1858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_1, ack => maxPool3D_CP_1610_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_update_start_
      -- CP-element group 30: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_sample_completed_
      -- 
    ra_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_673_inst_ack_0, ack => maxPool3D_CP_1610_elements(30)); -- 
    cr_1871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(30), ack => RPIPE_maxpool_input_pipe_673_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_673_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Sample/$entry
      -- 
    ca_1872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_673_inst_ack_1, ack => maxPool3D_CP_1610_elements(31)); -- 
    rr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(31), ack => type_cast_677_inst_req_0); -- 
    rr_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(31), ack => RPIPE_maxpool_input_pipe_685_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Sample/ra
      -- 
    ra_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_0, ack => maxPool3D_CP_1610_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	50 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_677_Update/$exit
      -- 
    ca_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_1, ack => maxPool3D_CP_1610_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_update_start_
      -- CP-element group 34: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_sample_completed_
      -- 
    ra_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_685_inst_ack_0, ack => maxPool3D_CP_1610_elements(34)); -- 
    cr_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(34), ack => RPIPE_maxpool_input_pipe_685_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_685_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Sample/rr
      -- 
    ca_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_685_inst_ack_1, ack => maxPool3D_CP_1610_elements(35)); -- 
    rr_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(35), ack => type_cast_689_inst_req_0); -- 
    rr_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(35), ack => RPIPE_maxpool_input_pipe_698_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Sample/ra
      -- 
    ra_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_0, ack => maxPool3D_CP_1610_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	50 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_689_Update/ca
      -- 
    ca_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_1, ack => maxPool3D_CP_1610_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_update_start_
      -- CP-element group 38: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Update/cr
      -- 
    ra_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_698_inst_ack_0, ack => maxPool3D_CP_1610_elements(38)); -- 
    cr_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(38), ack => RPIPE_maxpool_input_pipe_698_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_698_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Sample/rr
      -- 
    ca_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_698_inst_ack_1, ack => maxPool3D_CP_1610_elements(39)); -- 
    rr_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(39), ack => type_cast_702_inst_req_0); -- 
    rr_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(39), ack => RPIPE_maxpool_input_pipe_710_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Sample/ra
      -- 
    ra_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_702_inst_ack_0, ack => maxPool3D_CP_1610_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_702_Update/ca
      -- 
    ca_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_702_inst_ack_1, ack => maxPool3D_CP_1610_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_update_start_
      -- CP-element group 42: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Update/cr
      -- 
    ra_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_710_inst_ack_0, ack => maxPool3D_CP_1610_elements(42)); -- 
    cr_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(42), ack => RPIPE_maxpool_input_pipe_710_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_710_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Sample/rr
      -- 
    ca_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_710_inst_ack_1, ack => maxPool3D_CP_1610_elements(43)); -- 
    rr_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(43), ack => type_cast_714_inst_req_0); -- 
    rr_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(43), ack => RPIPE_maxpool_input_pipe_723_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Sample/ra
      -- 
    ra_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_0, ack => maxPool3D_CP_1610_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_714_Update/ca
      -- 
    ca_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_1, ack => maxPool3D_CP_1610_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_update_start_
      -- CP-element group 46: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Update/cr
      -- 
    ra_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_723_inst_ack_0, ack => maxPool3D_CP_1610_elements(46)); -- 
    cr_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(46), ack => RPIPE_maxpool_input_pipe_723_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/RPIPE_maxpool_input_pipe_723_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Sample/rr
      -- 
    ca_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_723_inst_ack_1, ack => maxPool3D_CP_1610_elements(47)); -- 
    rr_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(47), ack => type_cast_727_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Sample/ra
      -- 
    ra_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => maxPool3D_CP_1610_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/type_cast_727_Update/ca
      -- 
    ca_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => maxPool3D_CP_1610_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	21 
    -- CP-element group 50: 	29 
    -- CP-element group 50: 	33 
    -- CP-element group 50: 	37 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	9 
    -- CP-element group 50: 	13 
    -- CP-element group 50: 	17 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733/$exit
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_586_to_assign_stmt_733__exit__
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754__entry__
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/$entry
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_update_start_
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Update/cr
      -- 
    rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(50), ack => type_cast_737_inst_req_0); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(50), ack => type_cast_737_inst_req_1); -- 
    maxPool3D_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(25) & maxPool3D_CP_1610_elements(21) & maxPool3D_CP_1610_elements(29) & maxPool3D_CP_1610_elements(33) & maxPool3D_CP_1610_elements(37) & maxPool3D_CP_1610_elements(41) & maxPool3D_CP_1610_elements(45) & maxPool3D_CP_1610_elements(49) & maxPool3D_CP_1610_elements(5) & maxPool3D_CP_1610_elements(9) & maxPool3D_CP_1610_elements(13) & maxPool3D_CP_1610_elements(17);
      gj_maxPool3D_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Sample/ra
      -- 
    ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_737_inst_ack_0, ack => maxPool3D_CP_1610_elements(51)); -- 
    -- CP-element group 52:  branch  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (13) 
      -- CP-element group 52: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754__exit__
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755__entry__
      -- CP-element group 52: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/$exit
      -- CP-element group 52: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_583/assign_stmt_738_to_assign_stmt_754/type_cast_737_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755_dead_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755_eval_test/$entry
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755_eval_test/$exit
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755_eval_test/branch_req
      -- CP-element group 52: 	 branch_block_stmt_583/R_cmp195_756_place
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755_if_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_583/if_stmt_755_else_link/$entry
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_737_inst_ack_1, ack => maxPool3D_CP_1610_elements(52)); -- 
    branch_req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(52), ack => if_stmt_755_branch_req_0); -- 
    -- CP-element group 53:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (18) 
      -- CP-element group 53: 	 branch_block_stmt_583/merge_stmt_761_PhiAck/$exit
      -- CP-element group 53: 	 branch_block_stmt_583/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_583/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_583/merge_stmt_761_PhiReqMerge
      -- CP-element group 53: 	 branch_block_stmt_583/merge_stmt_761_PhiAck/dummy
      -- CP-element group 53: 	 branch_block_stmt_583/merge_stmt_761__exit__
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806__entry__
      -- CP-element group 53: 	 branch_block_stmt_583/merge_stmt_761_PhiAck/$entry
      -- CP-element group 53: 	 branch_block_stmt_583/if_stmt_755_if_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_583/if_stmt_755_if_link/if_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_583/entry_bbx_xnph
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/$entry
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_update_start_
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Update/cr
      -- 
    if_choice_transition_2028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_755_branch_ack_1, ack => maxPool3D_CP_1610_elements(53)); -- 
    rr_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(53), ack => type_cast_792_inst_req_0); -- 
    cr_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(53), ack => type_cast_792_inst_req_1); -- 
    -- CP-element group 54:  transition  place  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	204 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_583/if_stmt_755_else_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_583/if_stmt_755_else_link/else_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_583/entry_forx_xend
      -- CP-element group 54: 	 branch_block_stmt_583/entry_forx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_583/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_755_branch_ack_0, ack => maxPool3D_CP_1610_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Sample/ra
      -- 
    ra_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_792_inst_ack_0, ack => maxPool3D_CP_1610_elements(55)); -- 
    -- CP-element group 56:  transition  place  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	198 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/phi_stmt_809/$entry
      -- CP-element group 56: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806__exit__
      -- CP-element group 56: 	 branch_block_stmt_583/bbx_xnph_forx_xbody
      -- CP-element group 56: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/$exit
      -- CP-element group 56: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_583/assign_stmt_766_to_assign_stmt_806/type_cast_792_Update/ca
      -- 
    ca_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_792_inst_ack_1, ack => maxPool3D_CP_1610_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	203 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Sample/cra
      -- 
    cra_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_818_call_ack_0, ack => maxPool3D_CP_1610_elements(57)); -- 
    -- CP-element group 58:  branch  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	203 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829__exit__
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830__entry__
      -- CP-element group 58: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/$exit
      -- CP-element group 58: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Update/cca
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_583/R_exitcond1_831_place
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_583/if_stmt_830_else_link/$entry
      -- 
    cca_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_818_call_ack_1, ack => maxPool3D_CP_1610_elements(58)); -- 
    branch_req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(58), ack => if_stmt_830_branch_req_0); -- 
    -- CP-element group 59:  merge  transition  place  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	204 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_583/merge_stmt_836__exit__
      -- CP-element group 59: 	 branch_block_stmt_583/forx_xendx_xloopexit_forx_xend
      -- CP-element group 59: 	 branch_block_stmt_583/if_stmt_830_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_583/if_stmt_830_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_583/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 59: 	 branch_block_stmt_583/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_583/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_583/merge_stmt_836_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_583/merge_stmt_836_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_583/merge_stmt_836_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_583/merge_stmt_836_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_583/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_583/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_830_branch_ack_1, ack => maxPool3D_CP_1610_elements(59)); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	199 
    -- CP-element group 60: 	200 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_583/if_stmt_830_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_583/if_stmt_830_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_830_branch_ack_0, ack => maxPool3D_CP_1610_elements(60)); -- 
    rr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(60), ack => type_cast_815_inst_req_0); -- 
    cr_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(60), ack => type_cast_815_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	204 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Sample/cra
      -- 
    cra_2102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_853_call_ack_0, ack => maxPool3D_CP_1610_elements(61)); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	204 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	65 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	67 
    -- CP-element group 62: 	68 
    -- CP-element group 62:  members (25) 
      -- CP-element group 62: 	 branch_block_stmt_583/call_stmt_853__exit__
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877__entry__
      -- CP-element group 62: 	 branch_block_stmt_583/call_stmt_853/$exit
      -- CP-element group 62: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Update/cca
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_update_start_
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_update_start_
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_update_start_
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Update/cr
      -- 
    cca_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_853_call_ack_1, ack => maxPool3D_CP_1610_elements(62)); -- 
    rr_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(62), ack => type_cast_857_inst_req_0); -- 
    cr_2123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(62), ack => type_cast_857_inst_req_1); -- 
    rr_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(62), ack => type_cast_861_inst_req_0); -- 
    cr_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(62), ack => type_cast_861_inst_req_1); -- 
    rr_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(62), ack => type_cast_865_inst_req_0); -- 
    cr_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(62), ack => type_cast_865_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Sample/ra
      -- 
    ra_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_0, ack => maxPool3D_CP_1610_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_857_Update/ca
      -- 
    ca_2124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_1, ack => maxPool3D_CP_1610_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	62 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Sample/ra
      -- 
    ra_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_0, ack => maxPool3D_CP_1610_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_861_Update/ca
      -- 
    ca_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_1, ack => maxPool3D_CP_1610_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	62 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Sample/ra
      -- 
    ra_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_865_inst_ack_0, ack => maxPool3D_CP_1610_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	62 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/type_cast_865_Update/ca
      -- 
    ca_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_865_inst_ack_1, ack => maxPool3D_CP_1610_elements(68)); -- 
    -- CP-element group 69:  join  transition  place  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	66 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (10) 
      -- CP-element group 69: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877__exit__
      -- CP-element group 69: 	 branch_block_stmt_583/forx_xend_whilex_xbody
      -- CP-element group 69: 	 branch_block_stmt_583/merge_stmt_879__exit__
      -- CP-element group 69: 	 branch_block_stmt_583/do_while_stmt_896__entry__
      -- CP-element group 69: 	 branch_block_stmt_583/assign_stmt_858_to_assign_stmt_877/$exit
      -- CP-element group 69: 	 branch_block_stmt_583/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_583/forx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_583/merge_stmt_879_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_583/merge_stmt_879_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_583/merge_stmt_879_PhiAck/$exit
      -- 
    maxPool3D_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(64) & maxPool3D_CP_1610_elements(66) & maxPool3D_CP_1610_elements(68);
      gj_maxPool3D_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  place  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	76 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_583/do_while_stmt_896/$entry
      -- CP-element group 70: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896__entry__
      -- 
    maxPool3D_CP_1610_elements(70) <= maxPool3D_CP_1610_elements(69);
    -- CP-element group 71:  merge  place  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	180 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896__exit__
      -- 
    -- Element group maxPool3D_CP_1610_elements(71) is bound as output of CP function.
    -- CP-element group 72:  merge  place  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_583/do_while_stmt_896/loop_back
      -- 
    -- Element group maxPool3D_CP_1610_elements(72) is bound as output of CP function.
    -- CP-element group 73:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	78 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	178 
    -- CP-element group 73: 	179 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_583/do_while_stmt_896/loop_taken/$entry
      -- CP-element group 73: 	 branch_block_stmt_583/do_while_stmt_896/loop_exit/$entry
      -- CP-element group 73: 	 branch_block_stmt_583/do_while_stmt_896/condition_done
      -- 
    maxPool3D_CP_1610_elements(73) <= maxPool3D_CP_1610_elements(78);
    -- CP-element group 74:  branch  place  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	177 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_583/do_while_stmt_896/loop_body_done
      -- 
    maxPool3D_CP_1610_elements(74) <= maxPool3D_CP_1610_elements(177);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	87 
    -- CP-element group 75: 	108 
    -- CP-element group 75: 	129 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/back_edge_to_loop_body
      -- 
    maxPool3D_CP_1610_elements(75) <= maxPool3D_CP_1610_elements(72);
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	70 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	89 
    -- CP-element group 76: 	110 
    -- CP-element group 76: 	131 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/first_time_through_loop_body
      -- 
    maxPool3D_CP_1610_elements(76) <= maxPool3D_CP_1610_elements(70);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	83 
    -- CP-element group 77: 	84 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	103 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	176 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/$entry
      -- CP-element group 77: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/loop_body_start
      -- 
    -- Element group maxPool3D_CP_1610_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	171 
    -- CP-element group 78: 	175 
    -- CP-element group 78: 	176 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	73 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/condition_evaluated
      -- 
    condition_evaluated_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(78), ack => do_while_stmt_896_branch_req_0); -- 
    maxPool3D_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(82) & maxPool3D_CP_1610_elements(171) & maxPool3D_CP_1610_elements(175) & maxPool3D_CP_1610_elements(176);
      gj_maxPool3D_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: 	102 
    -- CP-element group 79: 	123 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	104 
    -- CP-element group 79: 	125 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/aggregated_phi_sample_req
      -- CP-element group 79: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_sample_start__ps
      -- 
    maxPool3D_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(83) & maxPool3D_CP_1610_elements(102) & maxPool3D_CP_1610_elements(123) & maxPool3D_CP_1610_elements(82);
      gj_maxPool3D_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	85 
    -- CP-element group 80: 	105 
    -- CP-element group 80: 	126 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	161 
    -- CP-element group 80: 	165 
    -- CP-element group 80: 	169 
    -- CP-element group 80: 	173 
    -- CP-element group 80: 	177 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80: 	102 
    -- CP-element group 80: 	123 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/aggregated_phi_sample_ack
      -- CP-element group 80: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_sample_completed_
      -- 
    maxPool3D_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(85) & maxPool3D_CP_1610_elements(105) & maxPool3D_CP_1610_elements(126);
      gj_maxPool3D_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	84 
    -- CP-element group 81: 	103 
    -- CP-element group 81: 	124 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	106 
    -- CP-element group 81: 	127 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/aggregated_phi_update_req
      -- CP-element group 81: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_update_start__ps
      -- 
    maxPool3D_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(84) & maxPool3D_CP_1610_elements(103) & maxPool3D_CP_1610_elements(124);
      gj_maxPool3D_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	86 
    -- CP-element group 82: 	107 
    -- CP-element group 82: 	128 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/aggregated_phi_update_ack
      -- 
    maxPool3D_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(86) & maxPool3D_CP_1610_elements(107) & maxPool3D_CP_1610_elements(128);
      gj_maxPool3D_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	171 
    -- CP-element group 83: 	175 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_sample_start_
      -- 
    maxPool3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(77) & maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(171) & maxPool3D_CP_1610_elements(175);
      gj_maxPool3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: 	154 
    -- CP-element group 84: 	174 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	81 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_update_start_
      -- 
    maxPool3D_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(77) & maxPool3D_CP_1610_elements(86) & maxPool3D_CP_1610_elements(154) & maxPool3D_CP_1610_elements(174);
      gj_maxPool3D_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	80 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	152 
    -- CP-element group 86: 	172 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(86) is bound as output of CP function.
    -- CP-element group 87:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	75 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_loopback_trigger
      -- 
    maxPool3D_CP_1610_elements(87) <= maxPool3D_CP_1610_elements(75);
    -- CP-element group 88:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_loopback_sample_req
      -- CP-element group 88: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_loopback_sample_req_ps
      -- 
    phi_stmt_898_loopback_sample_req_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_898_loopback_sample_req_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(88), ack => phi_stmt_898_req_0); -- 
    -- Element group maxPool3D_CP_1610_elements(88) is bound as output of CP function.
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	76 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_entry_trigger
      -- 
    maxPool3D_CP_1610_elements(89) <= maxPool3D_CP_1610_elements(76);
    -- CP-element group 90:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_entry_sample_req
      -- CP-element group 90: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_entry_sample_req_ps
      -- 
    phi_stmt_898_entry_sample_req_2185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_898_entry_sample_req_2185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(90), ack => phi_stmt_898_req_1); -- 
    -- Element group maxPool3D_CP_1610_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_phi_mux_ack
      -- CP-element group 91: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_898_phi_mux_ack_ps
      -- 
    phi_stmt_898_phi_mux_ack_2188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_898_ack_0, ack => maxPool3D_CP_1610_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_update_start__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Sample/rr
      -- 
    rr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(94), ack => type_cast_901_inst_req_0); -- 
    maxPool3D_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(92) & maxPool3D_CP_1610_elements(96);
      gj_maxPool3D_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_update_start_
      -- CP-element group 95: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Update/cr
      -- 
    cr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(95), ack => type_cast_901_inst_req_1); -- 
    maxPool3D_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(93) & maxPool3D_CP_1610_elements(97);
      gj_maxPool3D_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Sample/ra
      -- 
    ra_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_901_inst_ack_0, ack => maxPool3D_CP_1610_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_update_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_901_Update/ca
      -- 
    ca_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_901_inst_ack_1, ack => maxPool3D_CP_1610_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_sample_start__ps
      -- CP-element group 98: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_sample_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_sample_completed_
      -- 
    -- Element group maxPool3D_CP_1610_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_update_start__ps
      -- CP-element group 99: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_update_start_
      -- 
    -- Element group maxPool3D_CP_1610_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_update_completed__ps
      -- 
    maxPool3D_CP_1610_elements(100) <= maxPool3D_CP_1610_elements(101);
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	100 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_rowx_x1_at_entry_902_update_completed_
      -- 
    -- Element group maxPool3D_CP_1610_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => maxPool3D_CP_1610_elements(99), ack => maxPool3D_CP_1610_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	80 
    -- CP-element group 102: 	163 
    -- CP-element group 102: 	167 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	79 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_sample_start_
      -- 
    maxPool3D_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(77) & maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(163) & maxPool3D_CP_1610_elements(167);
      gj_maxPool3D_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	77 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	107 
    -- CP-element group 103: 	150 
    -- CP-element group 103: 	166 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	81 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_update_start_
      -- 
    maxPool3D_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(77) & maxPool3D_CP_1610_elements(107) & maxPool3D_CP_1610_elements(150) & maxPool3D_CP_1610_elements(166);
      gj_maxPool3D_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	79 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_sample_start__ps
      -- 
    maxPool3D_CP_1610_elements(104) <= maxPool3D_CP_1610_elements(79);
    -- CP-element group 105:  join  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	80 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	81 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_update_start__ps
      -- 
    maxPool3D_CP_1610_elements(106) <= maxPool3D_CP_1610_elements(81);
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	82 
    -- CP-element group 107: 	148 
    -- CP-element group 107: 	164 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	103 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	75 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_loopback_trigger
      -- 
    maxPool3D_CP_1610_elements(108) <= maxPool3D_CP_1610_elements(75);
    -- CP-element group 109:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_loopback_sample_req
      -- CP-element group 109: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_loopback_sample_req_ps
      -- 
    phi_stmt_903_loopback_sample_req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_903_loopback_sample_req_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(109), ack => phi_stmt_903_req_0); -- 
    -- Element group maxPool3D_CP_1610_elements(109) is bound as output of CP function.
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_entry_trigger
      -- 
    maxPool3D_CP_1610_elements(110) <= maxPool3D_CP_1610_elements(76);
    -- CP-element group 111:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_entry_sample_req
      -- CP-element group 111: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_entry_sample_req_ps
      -- 
    phi_stmt_903_entry_sample_req_2229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_903_entry_sample_req_2229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(111), ack => phi_stmt_903_req_1); -- 
    -- Element group maxPool3D_CP_1610_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_phi_mux_ack
      -- CP-element group 112: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_903_phi_mux_ack_ps
      -- 
    phi_stmt_903_phi_mux_ack_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_903_ack_0, ack => maxPool3D_CP_1610_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_update_start__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_sample_start_
      -- 
    rr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(115), ack => type_cast_906_inst_req_0); -- 
    maxPool3D_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(113) & maxPool3D_CP_1610_elements(117);
      gj_maxPool3D_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_update_start_
      -- 
    cr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(116), ack => type_cast_906_inst_req_1); -- 
    maxPool3D_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(114) & maxPool3D_CP_1610_elements(118);
      gj_maxPool3D_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_sample_completed__ps
      -- 
    ra_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_0, ack => maxPool3D_CP_1610_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_906_update_completed__ps
      -- 
    ca_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_1, ack => maxPool3D_CP_1610_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_sample_start__ps
      -- CP-element group 119: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_sample_completed__ps
      -- CP-element group 119: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_sample_completed_
      -- 
    -- Element group maxPool3D_CP_1610_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_update_start__ps
      -- CP-element group 120: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_update_start_
      -- 
    -- Element group maxPool3D_CP_1610_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_update_completed__ps
      -- 
    maxPool3D_CP_1610_elements(121) <= maxPool3D_CP_1610_elements(122);
    -- CP-element group 122:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	121 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_colx_x1_at_entry_907_update_completed_
      -- 
    -- Element group maxPool3D_CP_1610_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => maxPool3D_CP_1610_elements(120), ack => maxPool3D_CP_1610_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	80 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	79 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_sample_start_
      -- 
    maxPool3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(77) & maxPool3D_CP_1610_elements(80);
      gj_maxPool3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	128 
    -- CP-element group 124: 	146 
    -- CP-element group 124: 	162 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	81 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_update_start_
      -- 
    maxPool3D_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(77) & maxPool3D_CP_1610_elements(128) & maxPool3D_CP_1610_elements(146) & maxPool3D_CP_1610_elements(162);
      gj_maxPool3D_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_sample_start__ps
      -- 
    maxPool3D_CP_1610_elements(125) <= maxPool3D_CP_1610_elements(79);
    -- CP-element group 126:  join  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	80 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(126) is bound as output of CP function.
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	81 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_update_start__ps
      -- 
    maxPool3D_CP_1610_elements(127) <= maxPool3D_CP_1610_elements(81);
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	82 
    -- CP-element group 128: 	144 
    -- CP-element group 128: 	160 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	124 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(128) is bound as output of CP function.
    -- CP-element group 129:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	75 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_loopback_trigger
      -- 
    maxPool3D_CP_1610_elements(129) <= maxPool3D_CP_1610_elements(75);
    -- CP-element group 130:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_loopback_sample_req_ps
      -- CP-element group 130: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_loopback_sample_req
      -- 
    phi_stmt_908_loopback_sample_req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_908_loopback_sample_req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(130), ack => phi_stmt_908_req_0); -- 
    -- Element group maxPool3D_CP_1610_elements(130) is bound as output of CP function.
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	76 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_entry_trigger
      -- 
    maxPool3D_CP_1610_elements(131) <= maxPool3D_CP_1610_elements(76);
    -- CP-element group 132:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_entry_sample_req_ps
      -- CP-element group 132: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_entry_sample_req
      -- 
    phi_stmt_908_entry_sample_req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_908_entry_sample_req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(132), ack => phi_stmt_908_req_1); -- 
    -- Element group maxPool3D_CP_1610_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_phi_mux_ack_ps
      -- CP-element group 133: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/phi_stmt_908_phi_mux_ack
      -- 
    phi_stmt_908_phi_mux_ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_908_ack_0, ack => maxPool3D_CP_1610_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_update_start__ps
      -- 
    -- Element group maxPool3D_CP_1610_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_sample_start_
      -- 
    rr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(136), ack => type_cast_911_inst_req_0); -- 
    maxPool3D_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(134) & maxPool3D_CP_1610_elements(138);
      gj_maxPool3D_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_update_start_
      -- 
    cr_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(137), ack => type_cast_911_inst_req_1); -- 
    maxPool3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(135) & maxPool3D_CP_1610_elements(139);
      gj_maxPool3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_sample_completed__ps
      -- 
    ra_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_911_inst_ack_0, ack => maxPool3D_CP_1610_elements(138)); -- 
    -- CP-element group 139:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_911_update_completed__ps
      -- 
    ca_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_911_inst_ack_1, ack => maxPool3D_CP_1610_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_sample_completed_
      -- 
    -- Element group maxPool3D_CP_1610_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_update_start_
      -- 
    -- Element group maxPool3D_CP_1610_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_update_completed__ps
      -- 
    maxPool3D_CP_1610_elements(142) <= maxPool3D_CP_1610_elements(143);
    -- CP-element group 143:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/R_chlx_x0_at_entry_912_update_completed_
      -- 
    -- Element group maxPool3D_CP_1610_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => maxPool3D_CP_1610_elements(141), ack => maxPool3D_CP_1610_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	128 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Sample/rr
      -- 
    rr_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(144), ack => type_cast_916_inst_req_0); -- 
    maxPool3D_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(128) & maxPool3D_CP_1610_elements(146);
      gj_maxPool3D_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	158 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_update_start_
      -- 
    cr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(145), ack => type_cast_916_inst_req_1); -- 
    maxPool3D_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(147) & maxPool3D_CP_1610_elements(158);
      gj_maxPool3D_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	124 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Sample/ra
      -- 
    ra_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => maxPool3D_CP_1610_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	156 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_916_update_completed_
      -- 
    ca_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => maxPool3D_CP_1610_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	107 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_sample_start_
      -- 
    rr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(148), ack => type_cast_920_inst_req_0); -- 
    maxPool3D_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(107) & maxPool3D_CP_1610_elements(150);
      gj_maxPool3D_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	158 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_update_start_
      -- 
    cr_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(149), ack => type_cast_920_inst_req_1); -- 
    maxPool3D_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(151) & maxPool3D_CP_1610_elements(158);
      gj_maxPool3D_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	103 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_sample_completed_
      -- 
    ra_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_920_inst_ack_0, ack => maxPool3D_CP_1610_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	156 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_920_update_completed_
      -- 
    ca_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_920_inst_ack_1, ack => maxPool3D_CP_1610_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	86 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Sample/rr
      -- CP-element group 152: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_sample_start_
      -- 
    rr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(152), ack => type_cast_924_inst_req_0); -- 
    maxPool3D_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(86) & maxPool3D_CP_1610_elements(154);
      gj_maxPool3D_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	158 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_update_start_
      -- 
    cr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(153), ack => type_cast_924_inst_req_1); -- 
    maxPool3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(155) & maxPool3D_CP_1610_elements(158);
      gj_maxPool3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	84 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_sample_completed_
      -- 
    ra_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_0, ack => maxPool3D_CP_1610_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_924_update_completed_
      -- 
    ca_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_1, ack => maxPool3D_CP_1610_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	147 
    -- CP-element group 156: 	151 
    -- CP-element group 156: 	155 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Sample/crr
      -- CP-element group 156: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_sample_start_
      -- 
    crr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(156), ack => call_stmt_987_call_req_0); -- 
    maxPool3D_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(147) & maxPool3D_CP_1610_elements(151) & maxPool3D_CP_1610_elements(155) & maxPool3D_CP_1610_elements(158);
      gj_maxPool3D_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Update/ccr
      -- CP-element group 157: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_update_start_
      -- 
    ccr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(157), ack => call_stmt_987_call_req_1); -- 
    maxPool3D_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool3D_CP_1610_elements(159);
      gj_maxPool3D_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	145 
    -- CP-element group 158: 	149 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Sample/cra
      -- CP-element group 158: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_sample_completed_
      -- 
    cra_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_987_call_ack_0, ack => maxPool3D_CP_1610_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	177 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_Update/cca
      -- CP-element group 159: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/call_stmt_987_update_completed_
      -- 
    cca_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_987_call_ack_1, ack => maxPool3D_CP_1610_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	128 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Sample/rr
      -- 
    rr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(160), ack => type_cast_1001_inst_req_0); -- 
    maxPool3D_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(128) & maxPool3D_CP_1610_elements(162);
      gj_maxPool3D_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	80 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	170 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_update_start_
      -- CP-element group 161: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Update/cr
      -- 
    cr_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(161), ack => type_cast_1001_inst_req_1); -- 
    maxPool3D_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(163) & maxPool3D_CP_1610_elements(170);
      gj_maxPool3D_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	124 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Sample/ra
      -- 
    ra_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1001_inst_ack_0, ack => maxPool3D_CP_1610_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	168 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	102 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1001_Update/ca
      -- 
    ca_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1001_inst_ack_1, ack => maxPool3D_CP_1610_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	107 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Sample/req
      -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(164), ack => W_colx_x1_1002_delayed_1_0_1003_inst_req_0); -- 
    maxPool3D_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(107) & maxPool3D_CP_1610_elements(166);
      gj_maxPool3D_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	80 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	170 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_update_start_
      -- CP-element group 165: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Update/req
      -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(165), ack => W_colx_x1_1002_delayed_1_0_1003_inst_req_1); -- 
    maxPool3D_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(167) & maxPool3D_CP_1610_elements(170);
      gj_maxPool3D_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	103 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Sample/ack
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1002_delayed_1_0_1003_inst_ack_0, ack => maxPool3D_CP_1610_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	102 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1005_Update/ack
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1002_delayed_1_0_1003_inst_ack_1, ack => maxPool3D_CP_1610_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	163 
    -- CP-element group 168: 	167 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_sample_start_
      -- 
    rr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(168), ack => type_cast_1025_inst_req_0); -- 
    maxPool3D_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(163) & maxPool3D_CP_1610_elements(167) & maxPool3D_CP_1610_elements(170);
      gj_maxPool3D_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	80 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Update/cr
      -- CP-element group 169: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_update_start_
      -- 
    cr_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(169), ack => type_cast_1025_inst_req_1); -- 
    maxPool3D_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(171);
      gj_maxPool3D_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	161 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_sample_completed_
      -- 
    ra_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_0, ack => maxPool3D_CP_1610_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	78 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	83 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/type_cast_1025_Update/ca
      -- 
    ca_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_1, ack => maxPool3D_CP_1610_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	86 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Sample/req
      -- CP-element group 172: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_sample_start_
      -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(172), ack => W_rowx_x1_1023_delayed_2_0_1027_inst_req_0); -- 
    maxPool3D_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(86) & maxPool3D_CP_1610_elements(174);
      gj_maxPool3D_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	80 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Update/req
      -- CP-element group 173: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_update_start_
      -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(173), ack => W_rowx_x1_1023_delayed_2_0_1027_inst_req_1); -- 
    maxPool3D_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(175);
      gj_maxPool3D_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	84 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Sample/ack
      -- CP-element group 174: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_sample_completed_
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1023_delayed_2_0_1027_inst_ack_0, ack => maxPool3D_CP_1610_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	78 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	83 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Update/ack
      -- CP-element group 175: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/assign_stmt_1029_update_completed_
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1023_delayed_2_0_1027_inst_ack_1, ack => maxPool3D_CP_1610_elements(175)); -- 
    -- CP-element group 176:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	77 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	78 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group maxPool3D_CP_1610_elements(176) is a control-delay.
    cp_element_176_delay: control_delay_element  generic map(name => " 176_delay", delay_value => 1)  port map(req => maxPool3D_CP_1610_elements(77), ack => maxPool3D_CP_1610_elements(176), clk => clk, reset =>reset);
    -- CP-element group 177:  join  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	80 
    -- CP-element group 177: 	159 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	74 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_583/do_while_stmt_896/do_while_stmt_896_loop_body/$exit
      -- 
    maxPool3D_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(80) & maxPool3D_CP_1610_elements(159);
      gj_maxPool3D_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	73 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_583/do_while_stmt_896/loop_exit/ack
      -- CP-element group 178: 	 branch_block_stmt_583/do_while_stmt_896/loop_exit/$exit
      -- 
    ack_2421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_896_branch_ack_0, ack => maxPool3D_CP_1610_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	73 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_583/do_while_stmt_896/loop_taken/ack
      -- CP-element group 179: 	 branch_block_stmt_583/do_while_stmt_896/loop_taken/$exit
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_896_branch_ack_1, ack => maxPool3D_CP_1610_elements(179)); -- 
    -- CP-element group 180:  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	71 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	1 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_583/do_while_stmt_896/$exit
      -- 
    maxPool3D_CP_1610_elements(180) <= maxPool3D_CP_1610_elements(71);
    -- CP-element group 181:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	1 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	184 
    -- CP-element group 181:  members (18) 
      -- CP-element group 181: 	 branch_block_stmt_583/if_stmt_1053_if_link/$exit
      -- CP-element group 181: 	 branch_block_stmt_583/if_stmt_1053_if_link/if_choice_transition
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/$entry
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_update_start_
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_583/merge_stmt_1057__exit__
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063__entry__
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_583/whilex_xbody_whilex_xend
      -- CP-element group 181: 	 branch_block_stmt_583/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 181: 	 branch_block_stmt_583/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 181: 	 branch_block_stmt_583/merge_stmt_1057_PhiReqMerge
      -- CP-element group 181: 	 branch_block_stmt_583/merge_stmt_1057_PhiAck/$entry
      -- CP-element group 181: 	 branch_block_stmt_583/merge_stmt_1057_PhiAck/$exit
      -- CP-element group 181: 	 branch_block_stmt_583/merge_stmt_1057_PhiAck/dummy
      -- 
    if_choice_transition_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1053_branch_ack_1, ack => maxPool3D_CP_1610_elements(181)); -- 
    cr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(181), ack => type_cast_1062_inst_req_1); -- 
    rr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(181), ack => type_cast_1062_inst_req_0); -- 
    -- CP-element group 182:  merge  transition  place  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	1 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_583/if_stmt_1053_else_link/$exit
      -- CP-element group 182: 	 branch_block_stmt_583/if_stmt_1053_else_link/else_choice_transition
      -- CP-element group 182: 	 branch_block_stmt_583/if_stmt_1053__exit__
      -- CP-element group 182: 	 branch_block_stmt_583/merge_stmt_1057__entry__
      -- CP-element group 182: 	 branch_block_stmt_583/merge_stmt_1057_dead_link/$entry
      -- 
    else_choice_transition_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1053_branch_ack_0, ack => maxPool3D_CP_1610_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Sample/$exit
      -- 
    ra_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_0, ack => maxPool3D_CP_1610_elements(183)); -- 
    -- CP-element group 184:  fork  transition  place  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	181 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	186 
    -- CP-element group 184: 	188 
    -- CP-element group 184:  members (16) 
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Sample/crr
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Update/ccr
      -- CP-element group 184: 	 branch_block_stmt_583/assign_stmt_1063/$exit
      -- CP-element group 184: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_583/assign_stmt_1063__exit__
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079__entry__
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_update_start_
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/$entry
      -- CP-element group 184: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_update_start_
      -- CP-element group 184: 	 branch_block_stmt_583/assign_stmt_1063/type_cast_1062_Update/$exit
      -- 
    ca_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_1, ack => maxPool3D_CP_1610_elements(184)); -- 
    crr_2472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(184), ack => call_stmt_1066_call_req_0); -- 
    ccr_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(184), ack => call_stmt_1066_call_req_1); -- 
    cr_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(184), ack => type_cast_1070_inst_req_1); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Sample/cra
      -- CP-element group 185: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_sample_completed_
      -- 
    cra_2473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1066_call_ack_0, ack => maxPool3D_CP_1610_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/call_stmt_1066_Update/cca
      -- CP-element group 186: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Sample/$entry
      -- 
    cca_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1066_call_ack_1, ack => maxPool3D_CP_1610_elements(186)); -- 
    rr_2486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(186), ack => type_cast_1070_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Sample/$exit
      -- 
    ra_2487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_0, ack => maxPool3D_CP_1610_elements(187)); -- 
    -- CP-element group 188:  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	184 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (6) 
      -- CP-element group 188: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Sample/req
      -- CP-element group 188: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/type_cast_1070_update_completed_
      -- 
    ca_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_1, ack => maxPool3D_CP_1610_elements(188)); -- 
    req_2500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(188), ack => WPIPE_elapsed_time_pipe_1077_inst_req_0); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_update_start_
      -- CP-element group 189: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Sample/ack
      -- CP-element group 189: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Update/req
      -- CP-element group 189: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Update/$entry
      -- 
    ack_2501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1077_inst_ack_0, ack => maxPool3D_CP_1610_elements(189)); -- 
    req_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(189), ack => WPIPE_elapsed_time_pipe_1077_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  place  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	197 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	193 
    -- CP-element group 190: 	194 
    -- CP-element group 190:  members (22) 
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Update/ccr
      -- CP-element group 190: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_update_start_
      -- CP-element group 190: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079__exit__
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100__entry__
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/$exit
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_update_start_
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/$entry
      -- CP-element group 190: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Update/ack
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_583/call_stmt_1066_to_assign_stmt_1079/WPIPE_elapsed_time_pipe_1077_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_update_start_
      -- CP-element group 190: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_sample_start_
      -- 
    ack_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1077_inst_ack_1, ack => maxPool3D_CP_1610_elements(190)); -- 
    rr_2517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(190), ack => type_cast_1083_inst_req_0); -- 
    ccr_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(190), ack => call_stmt_1100_call_req_1); -- 
    cr_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(190), ack => type_cast_1083_inst_req_1); -- 
    cr_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(190), ack => type_cast_1087_inst_req_1); -- 
    rr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(190), ack => type_cast_1087_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_sample_completed_
      -- 
    ra_2518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_0, ack => maxPool3D_CP_1610_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1083_Update/ca
      -- 
    ca_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_1, ack => maxPool3D_CP_1610_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_sample_completed_
      -- 
    ra_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_0, ack => maxPool3D_CP_1610_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/type_cast_1087_update_completed_
      -- 
    ca_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_1, ack => maxPool3D_CP_1610_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Sample/crr
      -- CP-element group 195: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Sample/$entry
      -- 
    crr_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(195), ack => call_stmt_1100_call_req_0); -- 
    maxPool3D_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(192) & maxPool3D_CP_1610_elements(194);
      gj_maxPool3D_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Sample/cra
      -- CP-element group 196: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Sample/$exit
      -- 
    cra_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1100_call_ack_0, ack => maxPool3D_CP_1610_elements(196)); -- 
    -- CP-element group 197:  transition  place  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	190 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (16) 
      -- CP-element group 197: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Update/cca
      -- CP-element group 197: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_update_completed_
      -- CP-element group 197: 	 $exit
      -- CP-element group 197: 	 branch_block_stmt_583/$exit
      -- CP-element group 197: 	 branch_block_stmt_583/branch_block_stmt_583__exit__
      -- CP-element group 197: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100__exit__
      -- CP-element group 197: 	 branch_block_stmt_583/return__
      -- CP-element group 197: 	 branch_block_stmt_583/merge_stmt_1102__exit__
      -- CP-element group 197: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/call_stmt_1100_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_583/assign_stmt_1084_to_call_stmt_1100/$exit
      -- CP-element group 197: 	 branch_block_stmt_583/return___PhiReq/$entry
      -- CP-element group 197: 	 branch_block_stmt_583/return___PhiReq/$exit
      -- CP-element group 197: 	 branch_block_stmt_583/merge_stmt_1102_PhiReqMerge
      -- CP-element group 197: 	 branch_block_stmt_583/merge_stmt_1102_PhiAck/$entry
      -- CP-element group 197: 	 branch_block_stmt_583/merge_stmt_1102_PhiAck/$exit
      -- CP-element group 197: 	 branch_block_stmt_583/merge_stmt_1102_PhiAck/dummy
      -- 
    cca_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1100_call_ack_1, ack => maxPool3D_CP_1610_elements(197)); -- 
    -- CP-element group 198:  transition  output  delay-element  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	56 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	202 
    -- CP-element group 198:  members (5) 
      -- CP-element group 198: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/phi_stmt_809/$exit
      -- CP-element group 198: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 198: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/$exit
      -- CP-element group 198: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_813_konst_delay_trans
      -- CP-element group 198: 	 branch_block_stmt_583/bbx_xnph_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_req
      -- 
    phi_stmt_809_req_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_809_req_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(198), ack => phi_stmt_809_req_0); -- 
    -- Element group maxPool3D_CP_1610_elements(198) is a control-delay.
    cp_element_198_delay: control_delay_element  generic map(name => " 198_delay", delay_value => 1)  port map(req => maxPool3D_CP_1610_elements(56), ack => maxPool3D_CP_1610_elements(198), clk => clk, reset =>reset);
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	60 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Sample/ra
      -- 
    ra_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_0, ack => maxPool3D_CP_1610_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	60 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (2) 
      -- CP-element group 200: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/Update/ca
      -- 
    ca_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_1, ack => maxPool3D_CP_1610_elements(200)); -- 
    -- CP-element group 201:  join  transition  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 201: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/$exit
      -- CP-element group 201: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/$exit
      -- CP-element group 201: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/$exit
      -- CP-element group 201: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_sources/type_cast_815/SplitProtocol/$exit
      -- CP-element group 201: 	 branch_block_stmt_583/forx_xbody_forx_xbody_PhiReq/phi_stmt_809/phi_stmt_809_req
      -- 
    phi_stmt_809_req_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_809_req_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(201), ack => phi_stmt_809_req_1); -- 
    maxPool3D_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_1610_elements(199) & maxPool3D_CP_1610_elements(200);
      gj_maxPool3D_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_1610_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  merge  transition  place  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	198 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_583/merge_stmt_808_PhiReqMerge
      -- CP-element group 202: 	 branch_block_stmt_583/merge_stmt_808_PhiAck/$entry
      -- 
    maxPool3D_CP_1610_elements(202) <= OrReduce(maxPool3D_CP_1610_elements(198) & maxPool3D_CP_1610_elements(201));
    -- CP-element group 203:  fork  transition  place  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	57 
    -- CP-element group 203: 	58 
    -- CP-element group 203:  members (11) 
      -- CP-element group 203: 	 branch_block_stmt_583/merge_stmt_808__exit__
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829__entry__
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/$entry
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_update_start_
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Sample/crr
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_583/call_stmt_818_to_assign_stmt_829/call_stmt_818_Update/ccr
      -- CP-element group 203: 	 branch_block_stmt_583/merge_stmt_808_PhiAck/$exit
      -- CP-element group 203: 	 branch_block_stmt_583/merge_stmt_808_PhiAck/phi_stmt_809_ack
      -- 
    phi_stmt_809_ack_2605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_809_ack_0, ack => maxPool3D_CP_1610_elements(203)); -- 
    crr_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(203), ack => call_stmt_818_call_req_0); -- 
    ccr_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(203), ack => call_stmt_818_call_req_1); -- 
    -- CP-element group 204:  merge  fork  transition  place  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	54 
    -- CP-element group 204: 	59 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	61 
    -- CP-element group 204: 	62 
    -- CP-element group 204:  members (17) 
      -- CP-element group 204: 	 branch_block_stmt_583/merge_stmt_838__exit__
      -- CP-element group 204: 	 branch_block_stmt_583/assign_stmt_845_to_assign_stmt_850__entry__
      -- CP-element group 204: 	 branch_block_stmt_583/assign_stmt_845_to_assign_stmt_850__exit__
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853__entry__
      -- CP-element group 204: 	 branch_block_stmt_583/assign_stmt_845_to_assign_stmt_850/$entry
      -- CP-element group 204: 	 branch_block_stmt_583/assign_stmt_845_to_assign_stmt_850/$exit
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/$entry
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_update_start_
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Sample/crr
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_583/call_stmt_853/call_stmt_853_Update/ccr
      -- CP-element group 204: 	 branch_block_stmt_583/merge_stmt_838_PhiReqMerge
      -- CP-element group 204: 	 branch_block_stmt_583/merge_stmt_838_PhiAck/$entry
      -- CP-element group 204: 	 branch_block_stmt_583/merge_stmt_838_PhiAck/$exit
      -- CP-element group 204: 	 branch_block_stmt_583/merge_stmt_838_PhiAck/dummy
      -- 
    crr_2101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(204), ack => call_stmt_853_call_req_0); -- 
    ccr_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_1610_elements(204), ack => call_stmt_853_call_req_1); -- 
    maxPool3D_CP_1610_elements(204) <= OrReduce(maxPool3D_CP_1610_elements(54) & maxPool3D_CP_1610_elements(59));
    maxPool3D_do_while_stmt_896_terminator_2426: loop_terminator -- 
      generic map (name => " maxPool3D_do_while_stmt_896_terminator_2426", max_iterations_in_flight =>15) 
      port map(loop_body_exit => maxPool3D_CP_1610_elements(74),loop_continue => maxPool3D_CP_1610_elements(179),loop_terminate => maxPool3D_CP_1610_elements(178),loop_back => maxPool3D_CP_1610_elements(72),loop_exit => maxPool3D_CP_1610_elements(71),clk => clk, reset => reset); -- 
    phi_stmt_898_phi_seq_2216_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_1610_elements(87);
      maxPool3D_CP_1610_elements(92)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_1610_elements(96);
      maxPool3D_CP_1610_elements(93)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_1610_elements(97);
      maxPool3D_CP_1610_elements(88) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_1610_elements(89);
      maxPool3D_CP_1610_elements(98)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_1610_elements(98);
      maxPool3D_CP_1610_elements(99)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_1610_elements(100);
      maxPool3D_CP_1610_elements(90) <= phi_mux_reqs(1);
      phi_stmt_898_phi_seq_2216 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_898_phi_seq_2216") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_1610_elements(79), 
          phi_sample_ack => maxPool3D_CP_1610_elements(85), 
          phi_update_req => maxPool3D_CP_1610_elements(81), 
          phi_update_ack => maxPool3D_CP_1610_elements(86), 
          phi_mux_ack => maxPool3D_CP_1610_elements(91), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_903_phi_seq_2260_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_1610_elements(108);
      maxPool3D_CP_1610_elements(113)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_1610_elements(117);
      maxPool3D_CP_1610_elements(114)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_1610_elements(118);
      maxPool3D_CP_1610_elements(109) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_1610_elements(110);
      maxPool3D_CP_1610_elements(119)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_1610_elements(119);
      maxPool3D_CP_1610_elements(120)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_1610_elements(121);
      maxPool3D_CP_1610_elements(111) <= phi_mux_reqs(1);
      phi_stmt_903_phi_seq_2260 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_903_phi_seq_2260") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_1610_elements(104), 
          phi_sample_ack => maxPool3D_CP_1610_elements(105), 
          phi_update_req => maxPool3D_CP_1610_elements(106), 
          phi_update_ack => maxPool3D_CP_1610_elements(107), 
          phi_mux_ack => maxPool3D_CP_1610_elements(112), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_908_phi_seq_2304_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_1610_elements(129);
      maxPool3D_CP_1610_elements(134)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_1610_elements(138);
      maxPool3D_CP_1610_elements(135)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_1610_elements(139);
      maxPool3D_CP_1610_elements(130) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_1610_elements(131);
      maxPool3D_CP_1610_elements(140)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_1610_elements(140);
      maxPool3D_CP_1610_elements(141)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_1610_elements(142);
      maxPool3D_CP_1610_elements(132) <= phi_mux_reqs(1);
      phi_stmt_908_phi_seq_2304 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_908_phi_seq_2304") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_1610_elements(125), 
          phi_sample_ack => maxPool3D_CP_1610_elements(126), 
          phi_update_req => maxPool3D_CP_1610_elements(127), 
          phi_update_ack => maxPool3D_CP_1610_elements(128), 
          phi_mux_ack => maxPool3D_CP_1610_elements(133), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2168_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= maxPool3D_CP_1610_elements(75);
        preds(1)  <= maxPool3D_CP_1610_elements(76);
        entry_tmerge_2168 : transition_merge -- 
          generic map(name => " entry_tmerge_2168")
          port map (preds => preds, symbol_out => maxPool3D_CP_1610_elements(77));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_1052_wire : std_logic_vector(0 downto 0);
    signal add101_877 : std_logic_vector(31 downto 0);
    signal add117_935 : std_logic_vector(31 downto 0);
    signal add119_945 : std_logic_vector(31 downto 0);
    signal add131_955 : std_logic_vector(31 downto 0);
    signal add134_965 : std_logic_vector(31 downto 0);
    signal add13_633 : std_logic_vector(15 downto 0);
    signal add141_970 : std_logic_vector(31 downto 0);
    signal add145_975 : std_logic_vector(31 downto 0);
    signal add148_980 : std_logic_vector(31 downto 0);
    signal add23_658 : std_logic_vector(15 downto 0);
    signal add33_683 : std_logic_vector(15 downto 0);
    signal add43_708 : std_logic_vector(31 downto 0);
    signal add53_733 : std_logic_vector(15 downto 0);
    signal add_608 : std_logic_vector(31 downto 0);
    signal call11_624 : std_logic_vector(7 downto 0);
    signal call149_987 : std_logic_vector(7 downto 0);
    signal call16_636 : std_logic_vector(7 downto 0);
    signal call179_1066 : std_logic_vector(63 downto 0);
    signal call21_649 : std_logic_vector(7 downto 0);
    signal call26_661 : std_logic_vector(7 downto 0);
    signal call2_599 : std_logic_vector(7 downto 0);
    signal call31_674 : std_logic_vector(7 downto 0);
    signal call36_686 : std_logic_vector(7 downto 0);
    signal call41_699 : std_logic_vector(7 downto 0);
    signal call46_711 : std_logic_vector(7 downto 0);
    signal call51_724 : std_logic_vector(7 downto 0);
    signal call6_611 : std_logic_vector(7 downto 0);
    signal call89_853 : std_logic_vector(63 downto 0);
    signal call_586 : std_logic_vector(7 downto 0);
    signal chlx_x0_908 : std_logic_vector(15 downto 0);
    signal chlx_x0_at_entry_890 : std_logic_vector(15 downto 0);
    signal chlx_x1_1017 : std_logic_vector(15 downto 0);
    signal cmp156_998 : std_logic_vector(0 downto 0);
    signal cmp164_1022 : std_logic_vector(0 downto 0);
    signal cmp174_1046 : std_logic_vector(0 downto 0);
    signal cmp195_754 : std_logic_vector(0 downto 0);
    signal colx_x1_1002_delayed_1_0_1005 : std_logic_vector(15 downto 0);
    signal colx_x1_903 : std_logic_vector(15 downto 0);
    signal colx_x1_at_entry_885 : std_logic_vector(15 downto 0);
    signal colx_x2_1041 : std_logic_vector(15 downto 0);
    signal conv100_862 : std_logic_vector(31 downto 0);
    signal conv107_917 : std_logic_vector(31 downto 0);
    signal conv111_921 : std_logic_vector(31 downto 0);
    signal conv113_866 : std_logic_vector(31 downto 0);
    signal conv115_925 : std_logic_vector(31 downto 0);
    signal conv12_628 : std_logic_vector(15 downto 0);
    signal conv180_1071 : std_logic_vector(63 downto 0);
    signal conv188_1084 : std_logic_vector(31 downto 0);
    signal conv191_1088 : std_logic_vector(31 downto 0);
    signal conv19_640 : std_logic_vector(15 downto 0);
    signal conv1_590 : std_logic_vector(31 downto 0);
    signal conv22_653 : std_logic_vector(15 downto 0);
    signal conv29_665 : std_logic_vector(15 downto 0);
    signal conv32_678 : std_logic_vector(15 downto 0);
    signal conv39_690 : std_logic_vector(31 downto 0);
    signal conv3_603 : std_logic_vector(31 downto 0);
    signal conv42_703 : std_logic_vector(31 downto 0);
    signal conv49_715 : std_logic_vector(15 downto 0);
    signal conv52_728 : std_logic_vector(15 downto 0);
    signal conv59_738 : std_logic_vector(31 downto 0);
    signal conv90_1063 : std_logic_vector(63 downto 0);
    signal conv98_858 : std_logic_vector(31 downto 0);
    signal conv9_615 : std_logic_vector(15 downto 0);
    signal exitcond1_829 : std_logic_vector(0 downto 0);
    signal iNsTr_14_793 : std_logic_vector(63 downto 0);
    signal iNsTr_20_809 : std_logic_vector(63 downto 0);
    signal inc151_993 : std_logic_vector(15 downto 0);
    signal inc159_1002 : std_logic_vector(15 downto 0);
    signal inc159x_xcolx_x1_1010 : std_logic_vector(15 downto 0);
    signal inc168_1026 : std_logic_vector(15 downto 0);
    signal inc168x_xrowx_x1_1034 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_824 : std_logic_vector(63 downto 0);
    signal mul116_930 : std_logic_vector(31 downto 0);
    signal mul118_940 : std_logic_vector(31 downto 0);
    signal mul130_950 : std_logic_vector(31 downto 0);
    signal mul132_872 : std_logic_vector(31 downto 0);
    signal mul189_1093 : std_logic_vector(31 downto 0);
    signal mul192_1098 : std_logic_vector(31 downto 0);
    signal mul62_748 : std_logic_vector(31 downto 0);
    signal mul86_850 : std_logic_vector(15 downto 0);
    signal mul_743 : std_logic_vector(31 downto 0);
    signal rowx_x1_1023_delayed_2_0_1029 : std_logic_vector(15 downto 0);
    signal rowx_x1_898 : std_logic_vector(15 downto 0);
    signal rowx_x1_at_entry_880 : std_logic_vector(15 downto 0);
    signal shl10_621 : std_logic_vector(15 downto 0);
    signal shl133_960 : std_logic_vector(31 downto 0);
    signal shl20_646 : std_logic_vector(15 downto 0);
    signal shl30_671 : std_logic_vector(15 downto 0);
    signal shl40_696 : std_logic_vector(31 downto 0);
    signal shl50_721 : std_logic_vector(15 downto 0);
    signal shl_596 : std_logic_vector(31 downto 0);
    signal shr79193_845 : std_logic_vector(15 downto 0);
    signal sub_1076 : std_logic_vector(63 downto 0);
    signal tmp198_771 : std_logic_vector(31 downto 0);
    signal tmp199_777 : std_logic_vector(31 downto 0);
    signal tmp199x_xop_789 : std_logic_vector(31 downto 0);
    signal tmp200_783 : std_logic_vector(0 downto 0);
    signal tmp203_806 : std_logic_vector(63 downto 0);
    signal tmp_766 : std_logic_vector(31 downto 0);
    signal type_cast_1014_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1038_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1061_wire : std_logic_vector(63 downto 0);
    signal type_cast_1069_wire : std_logic_vector(63 downto 0);
    signal type_cast_594_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_619_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_669_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_694_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_752_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_787_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_797_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_804_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_813_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_815_wire : std_logic_vector(63 downto 0);
    signal type_cast_822_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_901_wire : std_logic_vector(15 downto 0);
    signal type_cast_906_wire : std_logic_vector(15 downto 0);
    signal type_cast_911_wire : std_logic_vector(15 downto 0);
    signal type_cast_991_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_whilex_xend_taken_1049 : std_logic_vector(0 downto 0);
    signal xx_xop_799 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    chlx_x0_at_entry_890 <= "0000000000000000";
    colx_x1_at_entry_885 <= "0000000000000000";
    rowx_x1_at_entry_880 <= "0000000000000000";
    type_cast_1014_wire_constant <= "0000000000000000";
    type_cast_1038_wire_constant <= "0000000000000000";
    type_cast_594_wire_constant <= "00000000000000000000000000001000";
    type_cast_619_wire_constant <= "0000000000001000";
    type_cast_644_wire_constant <= "0000000000001000";
    type_cast_669_wire_constant <= "0000000000001000";
    type_cast_694_wire_constant <= "00000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000001000";
    type_cast_752_wire_constant <= "00000000000000000000000000001111";
    type_cast_775_wire_constant <= "00000000000000000000000000000100";
    type_cast_781_wire_constant <= "00000000000000000000000000000001";
    type_cast_787_wire_constant <= "11111111111111111111111111111111";
    type_cast_797_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_804_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_813_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_822_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_843_wire_constant <= "0000000000000100";
    type_cast_870_wire_constant <= "00000000000000000000000000000001";
    type_cast_991_wire_constant <= "0000000000000001";
    phi_stmt_809: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_813_wire_constant & type_cast_815_wire;
      req <= phi_stmt_809_req_0 & phi_stmt_809_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_809",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_809_ack_0,
          idata => idata,
          odata => iNsTr_20_809,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_809
    phi_stmt_898: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_901_wire & rowx_x1_at_entry_880;
      req <= phi_stmt_898_req_0 & phi_stmt_898_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_898",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_898_ack_0,
          idata => idata,
          odata => rowx_x1_898,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_898
    phi_stmt_903: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_906_wire & colx_x1_at_entry_885;
      req <= phi_stmt_903_req_0 & phi_stmt_903_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_903",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_903_ack_0,
          idata => idata,
          odata => colx_x1_903,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_903
    phi_stmt_908: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_911_wire & chlx_x0_at_entry_890;
      req <= phi_stmt_908_req_0 & phi_stmt_908_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_908",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_908_ack_0,
          idata => idata,
          odata => chlx_x0_908,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_908
    -- flow-through select operator MUX_1016_inst
    chlx_x1_1017 <= type_cast_1014_wire_constant when (cmp156_998(0) /=  '0') else inc151_993;
    -- flow-through select operator MUX_1040_inst
    colx_x2_1041 <= type_cast_1038_wire_constant when (cmp164_1022(0) /=  '0') else inc159x_xcolx_x1_1010;
    -- flow-through select operator MUX_805_inst
    tmp203_806 <= xx_xop_799 when (tmp200_783(0) /=  '0') else type_cast_804_wire_constant;
    W_colx_x1_1002_delayed_1_0_1003_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_colx_x1_1002_delayed_1_0_1003_inst_req_0;
      W_colx_x1_1002_delayed_1_0_1003_inst_ack_0<= wack(0);
      rreq(0) <= W_colx_x1_1002_delayed_1_0_1003_inst_req_1;
      W_colx_x1_1002_delayed_1_0_1003_inst_ack_1<= rack(0);
      W_colx_x1_1002_delayed_1_0_1003_inst : InterlockBuffer generic map ( -- 
        name => "W_colx_x1_1002_delayed_1_0_1003_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_903,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => colx_x1_1002_delayed_1_0_1005,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rowx_x1_1023_delayed_2_0_1027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rowx_x1_1023_delayed_2_0_1027_inst_req_0;
      W_rowx_x1_1023_delayed_2_0_1027_inst_ack_0<= wack(0);
      rreq(0) <= W_rowx_x1_1023_delayed_2_0_1027_inst_req_1;
      W_rowx_x1_1023_delayed_2_0_1027_inst_ack_1<= rack(0);
      W_rowx_x1_1023_delayed_2_0_1027_inst : InterlockBuffer generic map ( -- 
        name => "W_rowx_x1_1023_delayed_2_0_1027_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowx_x1_1023_delayed_2_0_1029,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_1047_inst
    process(cmp174_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp174_1046(0 downto 0);
      whilex_xbody_whilex_xend_taken_1049 <= tmp_var; -- 
    end process;
    type_cast_1001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1001_inst_req_0;
      type_cast_1001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1001_inst_req_1;
      type_cast_1001_inst_ack_1<= rack(0);
      type_cast_1001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1001_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp156_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc159_1002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1025_inst_req_0;
      type_cast_1025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1025_inst_req_1;
      type_cast_1025_inst_ack_1<= rack(0);
      type_cast_1025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1025_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp164_1022,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc168_1026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1062_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1062_inst_req_0;
      type_cast_1062_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1062_inst_req_1;
      type_cast_1062_inst_ack_1<= rack(0);
      type_cast_1062_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1062_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1061_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1063,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1070_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1070_inst_req_0;
      type_cast_1070_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1070_inst_req_1;
      type_cast_1070_inst_ack_1<= rack(0);
      type_cast_1070_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1070_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1069_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv180_1071,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1083_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1083_inst_req_0;
      type_cast_1083_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1083_inst_req_1;
      type_cast_1083_inst_ack_1<= rack(0);
      type_cast_1083_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1083_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1087_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1087_inst_req_0;
      type_cast_1087_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1087_inst_req_1;
      type_cast_1087_inst_ack_1<= rack(0);
      type_cast_1087_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1087_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_1088,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_589_inst_req_0;
      type_cast_589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_589_inst_req_1;
      type_cast_589_inst_ack_1<= rack(0);
      type_cast_589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_602_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_602_inst_req_0;
      type_cast_602_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_602_inst_req_1;
      type_cast_602_inst_ack_1<= rack(0);
      type_cast_602_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_602_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_603,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_614_inst_req_0;
      type_cast_614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_614_inst_req_1;
      type_cast_614_inst_ack_1<= rack(0);
      type_cast_614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_627_inst_req_0;
      type_cast_627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_627_inst_req_1;
      type_cast_627_inst_ack_1<= rack(0);
      type_cast_627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_624,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_639_inst_req_0;
      type_cast_639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_639_inst_req_1;
      type_cast_639_inst_ack_1<= rack(0);
      type_cast_639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_652_inst_req_0;
      type_cast_652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_652_inst_req_1;
      type_cast_652_inst_ack_1<= rack(0);
      type_cast_652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_664_inst_req_0;
      type_cast_664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_664_inst_req_1;
      type_cast_664_inst_ack_1<= rack(0);
      type_cast_664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_677_inst_req_0;
      type_cast_677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_677_inst_req_1;
      type_cast_677_inst_ack_1<= rack(0);
      type_cast_677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_674,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_689_inst_req_0;
      type_cast_689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_689_inst_req_1;
      type_cast_689_inst_ack_1<= rack(0);
      type_cast_689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_702_inst_req_0;
      type_cast_702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_702_inst_req_1;
      type_cast_702_inst_ack_1<= rack(0);
      type_cast_702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_714_inst_req_0;
      type_cast_714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_714_inst_req_1;
      type_cast_714_inst_ack_1<= rack(0);
      type_cast_714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_737_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_737_inst_req_0;
      type_cast_737_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_737_inst_req_1;
      type_cast_737_inst_ack_1<= rack(0);
      type_cast_737_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_737_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_792_inst_req_0;
      type_cast_792_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_792_inst_req_1;
      type_cast_792_inst_ack_1<= rack(0);
      type_cast_792_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_792_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp199x_xop_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_793,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_815_inst_req_0;
      type_cast_815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_815_inst_req_1;
      type_cast_815_inst_ack_1<= rack(0);
      type_cast_815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_815_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_857_inst_req_0;
      type_cast_857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_857_inst_req_1;
      type_cast_857_inst_ack_1<= rack(0);
      type_cast_857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr79193_845,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_861_inst_req_0;
      type_cast_861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_861_inst_req_1;
      type_cast_861_inst_ack_1<= rack(0);
      type_cast_861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul86_850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_865_inst_req_0;
      type_cast_865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_865_inst_req_1;
      type_cast_865_inst_ack_1<= rack(0);
      type_cast_865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_901_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_901_inst_req_0;
      type_cast_901_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_901_inst_req_1;
      type_cast_901_inst_ack_1<= rack(0);
      type_cast_901_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_901_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc168x_xrowx_x1_1034,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_901_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_906_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_906_inst_req_0;
      type_cast_906_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_906_inst_req_1;
      type_cast_906_inst_ack_1<= rack(0);
      type_cast_906_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_906_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x2_1041,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_906_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_911_inst_req_0;
      type_cast_911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_911_inst_req_1;
      type_cast_911_inst_ack_1<= rack(0);
      type_cast_911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_911_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x1_1017,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_911_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x0_908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_917,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_920_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_920_inst_req_0;
      type_cast_920_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_920_inst_req_1;
      type_cast_920_inst_ack_1<= rack(0);
      type_cast_920_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_920_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_903,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_921,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_924_inst_req_0;
      type_cast_924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_924_inst_req_1;
      type_cast_924_inst_ack_1<= rack(0);
      type_cast_924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_896_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1052_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_896_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_896_branch_req_0,
          ack0 => do_while_stmt_896_branch_ack_0,
          ack1 => do_while_stmt_896_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1053_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_1049;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1053_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1053_branch_req_0,
          ack0 => if_stmt_1053_branch_ack_0,
          ack1 => if_stmt_1053_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_755_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp195_754;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_755_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_755_branch_req_0,
          ack0 => if_stmt_755_branch_ack_0,
          ack1 => if_stmt_755_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_830_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_829;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_830_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_830_branch_req_0,
          ack0 => if_stmt_830_branch_ack_0,
          ack1 => if_stmt_830_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1009_inst
    process(inc159_1002, colx_x1_1002_delayed_1_0_1005) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc159_1002, colx_x1_1002_delayed_1_0_1005, tmp_var);
      inc159x_xcolx_x1_1010 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1033_inst
    process(inc168_1026, rowx_x1_1023_delayed_2_0_1029) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc168_1026, rowx_x1_1023_delayed_2_0_1029, tmp_var);
      inc168x_xrowx_x1_1034 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_992_inst
    process(chlx_x0_908) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chlx_x0_908, type_cast_991_wire_constant, tmp_var);
      inc151_993 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_788_inst
    process(tmp199_777) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp199_777, type_cast_787_wire_constant, tmp_var);
      tmp199x_xop_789 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_876_inst
    process(conv100_862, conv98_858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv100_862, conv98_858, tmp_var);
      add101_877 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_934_inst
    process(conv111_921, mul116_930) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv111_921, mul116_930, tmp_var);
      add117_935 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_944_inst
    process(mul118_940, conv107_917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul118_940, conv107_917, tmp_var);
      add119_945 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_954_inst
    process(conv111_921, mul130_950) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv111_921, mul130_950, tmp_var);
      add131_955 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_964_inst
    process(shl133_960, conv107_917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl133_960, conv107_917, tmp_var);
      add134_965 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_969_inst
    process(add134_965, conv98_858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add134_965, conv98_858, tmp_var);
      add141_970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_974_inst
    process(add134_965, conv100_862) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add134_965, conv100_862, tmp_var);
      add145_975 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_979_inst
    process(add101_877, add134_965) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add101_877, add134_965, tmp_var);
      add148_980 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_798_inst
    process(iNsTr_14_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_14_793, type_cast_797_wire_constant, tmp_var);
      xx_xop_799 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_823_inst
    process(iNsTr_20_809) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_20_809, type_cast_822_wire_constant, tmp_var);
      indvarx_xnext_824 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1021_inst
    process(inc159x_xcolx_x1_1010, add33_683) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc159x_xcolx_x1_1010, add33_683, tmp_var);
      cmp164_1022 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1045_inst
    process(inc168x_xrowx_x1_1034, add13_633) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc168x_xrowx_x1_1034, add13_633, tmp_var);
      cmp174_1046 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_997_inst
    process(inc151_993, shr79193_845) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc151_993, shr79193_845, tmp_var);
      cmp156_998 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_828_inst
    process(indvarx_xnext_824, tmp203_806) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_824, tmp203_806, tmp_var);
      exitcond1_829 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_844_inst
    process(add53_733) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add53_733, type_cast_843_wire_constant, tmp_var);
      shr79193_845 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_776_inst
    process(tmp198_771) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp198_771, type_cast_775_wire_constant, tmp_var);
      tmp199_777 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_849_inst
    process(shr79193_845, add23_658) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(shr79193_845, add23_658, tmp_var);
      mul86_850 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1092_inst
    process(conv113_866, conv188_1084) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv113_866, conv188_1084, tmp_var);
      mul189_1093 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1097_inst
    process(mul189_1093, conv191_1088) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul189_1093, conv191_1088, tmp_var);
      mul192_1098 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_742_inst
    process(conv59_738, add_608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv59_738, add_608, tmp_var);
      mul_743 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_747_inst
    process(mul_743, add43_708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_743, add43_708, tmp_var);
      mul62_748 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_765_inst
    process(add_608, add43_708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_608, add43_708, tmp_var);
      tmp_766 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_770_inst
    process(tmp_766, conv59_738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_766, conv59_738, tmp_var);
      tmp198_771 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_929_inst
    process(conv115_925, conv113_866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv115_925, conv113_866, tmp_var);
      mul116_930 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_939_inst
    process(add117_935, conv98_858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add117_935, conv98_858, tmp_var);
      mul118_940 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_949_inst
    process(conv115_925, conv59_738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv115_925, conv59_738, tmp_var);
      mul130_950 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_959_inst
    process(mul132_872, add131_955) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul132_872, add131_955, tmp_var);
      shl133_960 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1052_inst
    process(cmp174_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp174_1046, tmp_var);
      NOT_u1_u1_1052_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_632_inst
    process(shl10_621, conv12_628) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_621, conv12_628, tmp_var);
      add13_633 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_657_inst
    process(shl20_646, conv22_653) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_646, conv22_653, tmp_var);
      add23_658 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_682_inst
    process(shl30_671, conv32_678) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_671, conv32_678, tmp_var);
      add33_683 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_732_inst
    process(shl50_721, conv52_728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_721, conv52_728, tmp_var);
      add53_733 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_607_inst
    process(shl_596, conv3_603) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_596, conv3_603, tmp_var);
      add_608 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_707_inst
    process(shl40_696, conv42_703) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_696, conv42_703, tmp_var);
      add43_708 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_620_inst
    process(conv9_615) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_615, type_cast_619_wire_constant, tmp_var);
      shl10_621 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_645_inst
    process(conv19_640) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_640, type_cast_644_wire_constant, tmp_var);
      shl20_646 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_670_inst
    process(conv29_665) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_665, type_cast_669_wire_constant, tmp_var);
      shl30_671 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_720_inst
    process(conv49_715) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_715, type_cast_719_wire_constant, tmp_var);
      shl50_721 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_595_inst
    process(conv1_590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_590, type_cast_594_wire_constant, tmp_var);
      shl_596 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_695_inst
    process(conv39_690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_690, type_cast_694_wire_constant, tmp_var);
      shl40_696 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_871_inst
    process(conv98_858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_858, type_cast_870_wire_constant, tmp_var);
      mul132_872 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1075_inst
    process(conv180_1071, conv90_1063) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv180_1071, conv90_1063, tmp_var);
      sub_1076 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_753_inst
    process(mul62_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul62_748, type_cast_752_wire_constant, tmp_var);
      cmp195_754 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_782_inst
    process(tmp199_777) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp199_777, type_cast_781_wire_constant, tmp_var);
      tmp200_783 <= tmp_var; --
    end process;
    -- unary operator type_cast_1061_inst
    process(call89_853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call89_853, tmp_var);
      type_cast_1061_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1069_inst
    process(call179_1066) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call179_1066, tmp_var);
      type_cast_1069_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_585_inst RPIPE_maxpool_input_pipe_598_inst RPIPE_maxpool_input_pipe_610_inst RPIPE_maxpool_input_pipe_623_inst RPIPE_maxpool_input_pipe_635_inst RPIPE_maxpool_input_pipe_648_inst RPIPE_maxpool_input_pipe_660_inst RPIPE_maxpool_input_pipe_673_inst RPIPE_maxpool_input_pipe_685_inst RPIPE_maxpool_input_pipe_698_inst RPIPE_maxpool_input_pipe_710_inst RPIPE_maxpool_input_pipe_723_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(95 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_585_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_598_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_610_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_623_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_635_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_648_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_660_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_673_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_685_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_698_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_710_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_723_inst_req_0;
      RPIPE_maxpool_input_pipe_585_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_598_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_610_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_623_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_635_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_648_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_660_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_673_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_685_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_698_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_710_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_723_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_585_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_598_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_610_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_623_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_635_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_648_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_660_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_673_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_685_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_698_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_710_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_723_inst_req_1;
      RPIPE_maxpool_input_pipe_585_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_598_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_610_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_623_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_635_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_648_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_660_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_673_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_685_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_698_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_710_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_723_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_586 <= data_out(95 downto 88);
      call2_599 <= data_out(87 downto 80);
      call6_611 <= data_out(79 downto 72);
      call11_624 <= data_out(71 downto 64);
      call16_636 <= data_out(63 downto 56);
      call21_649 <= data_out(55 downto 48);
      call26_661 <= data_out(47 downto 40);
      call31_674 <= data_out(39 downto 32);
      call36_686 <= data_out(31 downto 24);
      call41_699 <= data_out(23 downto 16);
      call46_711 <= data_out(15 downto 8);
      call51_724 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1077_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1077_inst_req_0;
      WPIPE_elapsed_time_pipe_1077_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1077_inst_req_1;
      WPIPE_elapsed_time_pipe_1077_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1076;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_853_call call_stmt_1066_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_853_call_req_0;
      reqL_unguarded(0) <= call_stmt_1066_call_req_0;
      call_stmt_853_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1066_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_853_call_req_1;
      reqR_unguarded(0) <= call_stmt_1066_call_req_1;
      call_stmt_853_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1066_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call89_853 <= data_out(127 downto 64);
      call179_1066 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1100_call 
    sendB_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1100_call_req_0;
      call_stmt_1100_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1100_call_req_1;
      call_stmt_1100_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_1_gI: SplitGuardInterface generic map(name => "sendB_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul192_1098;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(31 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_818_call 
    fill_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_818_call_req_0;
      call_stmt_818_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_818_call_req_1;
      call_stmt_818_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_T_call_group_2_gI: SplitGuardInterface generic map(name => "fill_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_20_809;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => fill_T_call_reqs(0),
          ackR => fill_T_call_acks(0),
          dataR => fill_T_call_data(63 downto 0),
          tagR => fill_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_T_return_acks(0), -- cross-over
          ackL => fill_T_return_reqs(0), -- cross-over
          tagL => fill_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_987_call 
    maxPool4_call_group_3: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 17);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_987_call_req_0;
      call_stmt_987_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_987_call_req_1;
      call_stmt_987_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      maxPool4_call_group_3_gI: SplitGuardInterface generic map(name => "maxPool4_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add119_945 & add134_965 & add141_970 & add145_975 & add148_980;
      call149_987 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 160,
        owidth => 160,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => maxPool4_call_reqs(0),
          ackR => maxPool4_call_acks(0),
          dataR => maxPool4_call_data(159 downto 0),
          tagR => maxPool4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => maxPool4_return_acks(0), -- cross-over
          ackL => maxPool4_return_reqs(0), -- cross-over
          dataL => maxPool4_return_data(7 downto 0),
          tagL => maxPool4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end maxPool3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    addr1 : in  std_logic_vector(31 downto 0);
    addr2 : in  std_logic_vector(31 downto 0);
    addr3 : in  std_logic_vector(31 downto 0);
    addr4 : in  std_logic_vector(31 downto 0);
    output : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool4;
architecture maxPool4_arch of maxPool4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 160)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal addr1_buffer :  std_logic_vector(31 downto 0);
  signal addr1_update_enable: Boolean;
  signal addr2_buffer :  std_logic_vector(31 downto 0);
  signal addr2_update_enable: Boolean;
  signal addr3_buffer :  std_logic_vector(31 downto 0);
  signal addr3_update_enable: Boolean;
  signal addr4_buffer :  std_logic_vector(31 downto 0);
  signal addr4_update_enable: Boolean;
  -- output port buffer signals
  signal output_buffer :  std_logic_vector(7 downto 0);
  signal output_update_enable: Boolean;
  signal maxPool4_CP_346_start: Boolean;
  signal maxPool4_CP_346_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_385_inst_ack_0 : boolean;
  signal type_cast_385_inst_req_0 : boolean;
  signal type_cast_385_inst_ack_1 : boolean;
  signal W_myptr5_366_delayed_8_0_366_inst_ack_0 : boolean;
  signal W_myptr5_366_delayed_8_0_366_inst_req_0 : boolean;
  signal type_cast_385_inst_req_1 : boolean;
  signal ptr_deref_370_store_0_ack_0 : boolean;
  signal addr_of_364_final_reg_req_0 : boolean;
  signal ptr_deref_370_store_0_req_0 : boolean;
  signal CONCAT_u32_u64_381_inst_ack_1 : boolean;
  signal addr_of_364_final_reg_ack_0 : boolean;
  signal CONCAT_u32_u64_381_inst_req_1 : boolean;
  signal CONCAT_u32_u64_381_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_381_inst_req_0 : boolean;
  signal addr_of_364_final_reg_ack_1 : boolean;
  signal ptr_deref_370_store_0_ack_1 : boolean;
  signal ptr_deref_119_load_0_req_0 : boolean;
  signal ptr_deref_119_load_0_ack_0 : boolean;
  signal ptr_deref_370_store_0_req_1 : boolean;
  signal W_myptr5_366_delayed_8_0_366_inst_ack_1 : boolean;
  signal addr_of_364_final_reg_req_1 : boolean;
  signal W_myptr5_366_delayed_8_0_366_inst_req_1 : boolean;
  signal array_obj_ref_93_index_offset_req_0 : boolean;
  signal array_obj_ref_93_index_offset_ack_0 : boolean;
  signal array_obj_ref_93_index_offset_req_1 : boolean;
  signal array_obj_ref_93_index_offset_ack_1 : boolean;
  signal addr_of_94_final_reg_req_0 : boolean;
  signal addr_of_94_final_reg_ack_0 : boolean;
  signal addr_of_94_final_reg_req_1 : boolean;
  signal addr_of_94_final_reg_ack_1 : boolean;
  signal array_obj_ref_100_index_offset_req_0 : boolean;
  signal array_obj_ref_100_index_offset_ack_0 : boolean;
  signal array_obj_ref_100_index_offset_req_1 : boolean;
  signal array_obj_ref_100_index_offset_ack_1 : boolean;
  signal addr_of_101_final_reg_req_0 : boolean;
  signal addr_of_101_final_reg_ack_0 : boolean;
  signal addr_of_101_final_reg_req_1 : boolean;
  signal addr_of_101_final_reg_ack_1 : boolean;
  signal array_obj_ref_107_index_offset_req_0 : boolean;
  signal array_obj_ref_107_index_offset_ack_0 : boolean;
  signal array_obj_ref_107_index_offset_req_1 : boolean;
  signal array_obj_ref_107_index_offset_ack_1 : boolean;
  signal addr_of_108_final_reg_req_0 : boolean;
  signal addr_of_108_final_reg_ack_0 : boolean;
  signal addr_of_108_final_reg_req_1 : boolean;
  signal addr_of_108_final_reg_ack_1 : boolean;
  signal array_obj_ref_114_index_offset_req_0 : boolean;
  signal array_obj_ref_114_index_offset_ack_0 : boolean;
  signal array_obj_ref_114_index_offset_req_1 : boolean;
  signal array_obj_ref_114_index_offset_ack_1 : boolean;
  signal addr_of_115_final_reg_req_0 : boolean;
  signal addr_of_115_final_reg_ack_0 : boolean;
  signal addr_of_115_final_reg_req_1 : boolean;
  signal addr_of_115_final_reg_ack_1 : boolean;
  signal ptr_deref_119_load_0_req_1 : boolean;
  signal ptr_deref_119_load_0_ack_1 : boolean;
  signal ptr_deref_123_load_0_req_0 : boolean;
  signal ptr_deref_123_load_0_ack_0 : boolean;
  signal ptr_deref_123_load_0_req_1 : boolean;
  signal ptr_deref_123_load_0_ack_1 : boolean;
  signal ptr_deref_127_load_0_req_0 : boolean;
  signal ptr_deref_127_load_0_ack_0 : boolean;
  signal ptr_deref_127_load_0_req_1 : boolean;
  signal ptr_deref_127_load_0_ack_1 : boolean;
  signal ptr_deref_131_load_0_req_0 : boolean;
  signal ptr_deref_131_load_0_ack_0 : boolean;
  signal ptr_deref_131_load_0_req_1 : boolean;
  signal ptr_deref_131_load_0_ack_1 : boolean;
  signal slice_136_inst_req_0 : boolean;
  signal slice_136_inst_ack_0 : boolean;
  signal slice_136_inst_req_1 : boolean;
  signal slice_136_inst_ack_1 : boolean;
  signal slice_140_inst_req_0 : boolean;
  signal slice_140_inst_ack_0 : boolean;
  signal slice_140_inst_req_1 : boolean;
  signal slice_140_inst_ack_1 : boolean;
  signal slice_144_inst_req_0 : boolean;
  signal slice_144_inst_ack_0 : boolean;
  signal slice_144_inst_req_1 : boolean;
  signal slice_144_inst_ack_1 : boolean;
  signal slice_148_inst_req_0 : boolean;
  signal slice_148_inst_ack_0 : boolean;
  signal slice_148_inst_req_1 : boolean;
  signal slice_148_inst_ack_1 : boolean;
  signal slice_152_inst_req_0 : boolean;
  signal slice_152_inst_ack_0 : boolean;
  signal slice_152_inst_req_1 : boolean;
  signal slice_152_inst_ack_1 : boolean;
  signal slice_156_inst_req_0 : boolean;
  signal slice_156_inst_ack_0 : boolean;
  signal slice_156_inst_req_1 : boolean;
  signal slice_156_inst_ack_1 : boolean;
  signal slice_160_inst_req_0 : boolean;
  signal slice_160_inst_ack_0 : boolean;
  signal slice_160_inst_req_1 : boolean;
  signal slice_160_inst_ack_1 : boolean;
  signal slice_164_inst_req_0 : boolean;
  signal slice_164_inst_ack_0 : boolean;
  signal slice_164_inst_req_1 : boolean;
  signal slice_164_inst_ack_1 : boolean;
  signal slice_168_inst_req_0 : boolean;
  signal slice_168_inst_ack_0 : boolean;
  signal slice_168_inst_req_1 : boolean;
  signal slice_168_inst_ack_1 : boolean;
  signal slice_172_inst_req_0 : boolean;
  signal slice_172_inst_ack_0 : boolean;
  signal slice_172_inst_req_1 : boolean;
  signal slice_172_inst_ack_1 : boolean;
  signal slice_176_inst_req_0 : boolean;
  signal slice_176_inst_ack_0 : boolean;
  signal slice_176_inst_req_1 : boolean;
  signal slice_176_inst_ack_1 : boolean;
  signal slice_180_inst_req_0 : boolean;
  signal slice_180_inst_ack_0 : boolean;
  signal slice_180_inst_req_1 : boolean;
  signal slice_180_inst_ack_1 : boolean;
  signal slice_184_inst_req_0 : boolean;
  signal slice_184_inst_ack_0 : boolean;
  signal slice_184_inst_req_1 : boolean;
  signal slice_184_inst_ack_1 : boolean;
  signal slice_188_inst_req_0 : boolean;
  signal slice_188_inst_ack_0 : boolean;
  signal slice_188_inst_req_1 : boolean;
  signal slice_188_inst_ack_1 : boolean;
  signal slice_192_inst_req_0 : boolean;
  signal slice_192_inst_ack_0 : boolean;
  signal slice_192_inst_req_1 : boolean;
  signal slice_192_inst_ack_1 : boolean;
  signal slice_196_inst_req_0 : boolean;
  signal slice_196_inst_ack_0 : boolean;
  signal slice_196_inst_req_1 : boolean;
  signal slice_196_inst_ack_1 : boolean;
  signal array_obj_ref_363_index_offset_req_0 : boolean;
  signal array_obj_ref_363_index_offset_ack_0 : boolean;
  signal array_obj_ref_363_index_offset_req_1 : boolean;
  signal array_obj_ref_363_index_offset_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool4_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 160) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= addr1;
  addr1_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(95 downto 64) <= addr2;
  addr2_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(127 downto 96) <= addr3;
  addr3_buffer <= in_buffer_data_out(127 downto 96);
  in_buffer_data_in(159 downto 128) <= addr4;
  addr4_buffer <= in_buffer_data_out(159 downto 128);
  in_buffer_data_in(tag_length + 159 downto 160) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 159 downto 160);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= addr_update_enable & addr1_update_enable & addr2_update_enable & addr3_update_enable & addr4_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool4_CP_346_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool4_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= output_buffer;
  output <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_346_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  output_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "output_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_output_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => output_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool4_CP_346_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_346_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool4_CP_346: Block -- control-path 
    signal maxPool4_CP_346_elements: BooleanArray(146 downto 0);
    -- 
  begin -- 
    maxPool4_CP_346_elements(0) <= maxPool4_CP_346_start;
    maxPool4_CP_346_symbol <= maxPool4_CP_346_elements(146);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	16 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	25 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	31 
    -- CP-element group 1: 	32 
    -- CP-element group 1: 	117 
    -- CP-element group 1: 	118 
    -- CP-element group 1: 	119 
    -- CP-element group 1:  members (66) 
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_resized_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_computed_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_resized_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_computed_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_resized_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_computed_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_resized_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_computed_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_resized_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_computed_1
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Sample/req
      -- 
    req_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_93_index_offset_req_0); -- 
    req_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_100_index_offset_req_0); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_107_index_offset_req_0); -- 
    req_526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_114_index_offset_req_0); -- 
    req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_363_index_offset_req_0); -- 
    maxPool4_CP_346_elements(1) <= maxPool4_CP_346_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	119 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	140 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_95_to_assign_stmt_386/addr_update_enable
      -- CP-element group 2: 	 assign_stmt_95_to_assign_stmt_386/addr_update_enable_out
      -- 
    maxPool4_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(119);
      gj_maxPool4_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	141 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_95_to_assign_stmt_386/addr1_update_enable
      -- CP-element group 3: 	 assign_stmt_95_to_assign_stmt_386/addr1_update_enable_out
      -- 
    maxPool4_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(11);
      gj_maxPool4_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	142 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_95_to_assign_stmt_386/addr2_update_enable
      -- CP-element group 4: 	 assign_stmt_95_to_assign_stmt_386/addr2_update_enable_out
      -- 
    maxPool4_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(18);
      gj_maxPool4_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	143 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_95_to_assign_stmt_386/addr3_update_enable
      -- CP-element group 5: 	 assign_stmt_95_to_assign_stmt_386/addr3_update_enable_out
      -- 
    maxPool4_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(25);
      gj_maxPool4_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	32 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	144 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_95_to_assign_stmt_386/addr4_update_enable
      -- CP-element group 6: 	 assign_stmt_95_to_assign_stmt_386/addr4_update_enable_out
      -- 
    maxPool4_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(32);
      gj_maxPool4_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	145 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	136 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_95_to_assign_stmt_386/output_update_enable
      -- CP-element group 7: 	 assign_stmt_95_to_assign_stmt_386/output_update_enable_in
      -- 
    maxPool4_CP_346_elements(7) <= maxPool4_CP_346_elements(145);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_sample_start_
      -- CP-element group 8: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_request/$entry
      -- CP-element group 8: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_request/req
      -- 
    req_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(8), ack => addr_of_94_final_reg_req_0); -- 
    maxPool4_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(12) & maxPool4_CP_346_elements(13);
      gj_maxPool4_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	38 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_update_start_
      -- CP-element group 9: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_complete/$entry
      -- CP-element group 9: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_complete/req
      -- 
    req_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(9), ack => addr_of_94_final_reg_req_1); -- 
    maxPool4_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(14) & maxPool4_CP_346_elements(38);
      gj_maxPool4_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_update_start
      -- CP-element group 10: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Update/$entry
      -- CP-element group 10: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Update/req
      -- 
    req_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(10), ack => array_obj_ref_93_index_offset_req_1); -- 
    maxPool4_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(12) & maxPool4_CP_346_elements(13);
      gj_maxPool4_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	139 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_sample_complete
      -- CP-element group 11: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Sample/ack
      -- 
    ack_389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_93_index_offset_ack_0, ack => maxPool4_CP_346_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_root_address_calculated
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_offset_calculated
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Update/$exit
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_final_index_sum_regn_Update/ack
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_base_plus_offset/$entry
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_base_plus_offset/$exit
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_93_base_plus_offset/sum_rename_ack
      -- 
    ack_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_93_index_offset_ack_1, ack => maxPool4_CP_346_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_sample_completed_
      -- CP-element group 13: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_request/$exit
      -- CP-element group 13: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_request/ack
      -- 
    ack_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_94_final_reg_ack_0, ack => maxPool4_CP_346_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (19) 
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_word_address_calculated
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_root_address_calculated
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_address_resized
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_addr_resize/$entry
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_addr_resize/$exit
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_addr_resize/base_resize_req
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_addr_resize/base_resize_ack
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_plus_offset/$entry
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_plus_offset/$exit
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_word_addrgen/$entry
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_word_addrgen/$exit
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_word_addrgen/root_register_req
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_word_addrgen/root_register_ack
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_update_completed_
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_complete/$exit
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/addr_of_94_complete/ack
      -- CP-element group 14: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_base_address_calculated
      -- 
    ack_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_94_final_reg_ack_1, ack => maxPool4_CP_346_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_sample_start_
      -- CP-element group 15: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_request/$entry
      -- CP-element group 15: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_request/req
      -- 
    req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(15), ack => addr_of_101_final_reg_req_0); -- 
    maxPool4_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(19) & maxPool4_CP_346_elements(20);
      gj_maxPool4_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	42 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_update_start_
      -- CP-element group 16: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_complete/$entry
      -- CP-element group 16: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_complete/req
      -- 
    req_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(16), ack => addr_of_101_final_reg_req_1); -- 
    maxPool4_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(21) & maxPool4_CP_346_elements(42);
      gj_maxPool4_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Update/req
      -- 
    req_439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(17), ack => array_obj_ref_100_index_offset_req_1); -- 
    maxPool4_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(19) & maxPool4_CP_346_elements(20);
      gj_maxPool4_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	139 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Sample/ack
      -- 
    ack_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_100_index_offset_ack_0, ack => maxPool4_CP_346_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (8) 
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_root_address_calculated
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_offset_calculated
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_base_plus_offset/$entry
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_base_plus_offset/$exit
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_100_base_plus_offset/sum_rename_ack
      -- 
    ack_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_100_index_offset_ack_1, ack => maxPool4_CP_346_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_sample_completed_
      -- CP-element group 20: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_request/$exit
      -- CP-element group 20: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_request/ack
      -- 
    ack_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_101_final_reg_ack_0, ack => maxPool4_CP_346_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	40 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_update_completed_
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_complete/$exit
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/addr_of_101_complete/ack
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_address_resized
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_word_addrgen/root_register_ack
      -- 
    ack_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_101_final_reg_ack_1, ack => maxPool4_CP_346_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_sample_start_
      -- CP-element group 22: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_request/$entry
      -- CP-element group 22: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_request/req
      -- 
    req_495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(22), ack => addr_of_108_final_reg_req_0); -- 
    maxPool4_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(26) & maxPool4_CP_346_elements(27);
      gj_maxPool4_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_update_start_
      -- CP-element group 23: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_complete/$entry
      -- CP-element group 23: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_complete/req
      -- 
    req_500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(23), ack => addr_of_108_final_reg_req_1); -- 
    maxPool4_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(28) & maxPool4_CP_346_elements(46);
      gj_maxPool4_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_update_start
      -- CP-element group 24: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Update/$entry
      -- CP-element group 24: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Update/req
      -- 
    req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(24), ack => array_obj_ref_107_index_offset_req_1); -- 
    maxPool4_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(26) & maxPool4_CP_346_elements(27);
      gj_maxPool4_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	1 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	139 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	5 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_sample_complete
      -- CP-element group 25: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Sample/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_107_index_offset_ack_0, ack => maxPool4_CP_346_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (8) 
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_offset_calculated
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Update/$exit
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_final_index_sum_regn_Update/ack
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_base_plus_offset/$exit
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_107_base_plus_offset/sum_rename_ack
      -- 
    ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_107_index_offset_ack_1, ack => maxPool4_CP_346_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	24 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_sample_completed_
      -- CP-element group 27: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_request/$exit
      -- CP-element group 27: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_request/ack
      -- 
    ack_496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_108_final_reg_ack_0, ack => maxPool4_CP_346_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	44 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28:  members (19) 
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_update_completed_
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_complete/$exit
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/addr_of_108_complete/ack
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_address_calculated
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_word_address_calculated
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_address_resized
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_addr_resize/$entry
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_addr_resize/$exit
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_addr_resize/base_resize_req
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_addr_resize/base_resize_ack
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_word_addrgen/$entry
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_word_addrgen/$exit
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_word_addrgen/root_register_req
      -- CP-element group 28: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_word_addrgen/root_register_ack
      -- 
    ack_501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_108_final_reg_ack_1, ack => maxPool4_CP_346_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	33 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	34 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_sample_start_
      -- CP-element group 29: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_request/$entry
      -- CP-element group 29: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_request/req
      -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(29), ack => addr_of_115_final_reg_req_0); -- 
    maxPool4_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(33) & maxPool4_CP_346_elements(34);
      gj_maxPool4_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	50 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_update_start_
      -- CP-element group 30: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_complete/$entry
      -- CP-element group 30: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_complete/req
      -- 
    req_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(30), ack => addr_of_115_final_reg_req_1); -- 
    maxPool4_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(35) & maxPool4_CP_346_elements(50);
      gj_maxPool4_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	1 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	34 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_update_start
      -- CP-element group 31: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Update/$entry
      -- CP-element group 31: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Update/req
      -- 
    req_531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(31), ack => array_obj_ref_114_index_offset_req_1); -- 
    maxPool4_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(33) & maxPool4_CP_346_elements(34);
      gj_maxPool4_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	1 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	139 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	6 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_sample_complete
      -- CP-element group 32: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Sample/ack
      -- 
    ack_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_114_index_offset_ack_0, ack => maxPool4_CP_346_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (8) 
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_root_address_calculated
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_offset_calculated
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_final_index_sum_regn_Update/ack
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_base_plus_offset/$entry
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_base_plus_offset/$exit
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_114_base_plus_offset/sum_rename_ack
      -- 
    ack_532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_114_index_offset_ack_1, ack => maxPool4_CP_346_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_sample_completed_
      -- CP-element group 34: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_request/$exit
      -- CP-element group 34: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_request/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_115_final_reg_ack_0, ack => maxPool4_CP_346_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	48 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	30 
    -- CP-element group 35:  members (19) 
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_root_address_calculated
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_update_completed_
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_complete/$exit
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/addr_of_115_complete/ack
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_address_calculated
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_word_address_calculated
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_address_resized
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_addr_resize/$entry
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_addr_resize/$exit
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_plus_offset/$entry
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_plus_offset/$exit
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_word_addrgen/$entry
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_word_addrgen/$exit
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_word_addrgen/root_register_req
      -- CP-element group 35: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_word_addrgen/root_register_ack
      -- 
    ack_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_115_final_reg_ack_1, ack => maxPool4_CP_346_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/word_access_start/$entry
      -- CP-element group 36: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/word_access_start/word_0/rr
      -- CP-element group 36: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_sample_start_
      -- 
    rr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(36), ack => ptr_deref_119_load_0_req_0); -- 
    maxPool4_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(14) & maxPool4_CP_346_elements(38);
      gj_maxPool4_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	66 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/$entry
      -- CP-element group 37: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_update_start_
      -- CP-element group 37: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/word_access_complete/$entry
      -- CP-element group 37: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/word_access_complete/word_0/cr
      -- 
    cr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(37), ack => ptr_deref_119_load_0_req_1); -- 
    maxPool4_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(54) & maxPool4_CP_346_elements(58) & maxPool4_CP_346_elements(62) & maxPool4_CP_346_elements(66);
      gj_maxPool4_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/word_access_start/$exit
      -- CP-element group 38: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Sample/word_access_start/word_0/ra
      -- CP-element group 38: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_sample_completed_
      -- 
    ra_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_119_load_0_ack_0, ack => maxPool4_CP_346_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	64 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/$exit
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_update_completed_
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/word_access_complete/$exit
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/ptr_deref_119_Merge/$entry
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/ptr_deref_119_Merge/$exit
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/ptr_deref_119_Merge/merge_req
      -- CP-element group 39: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_119_Update/ptr_deref_119_Merge/merge_ack
      -- 
    ca_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_119_load_0_ack_1, ack => maxPool4_CP_346_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	21 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_sample_start_
      -- CP-element group 40: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/word_access_start/$entry
      -- CP-element group 40: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/word_access_start/word_0/rr
      -- 
    rr_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(40), ack => ptr_deref_123_load_0_req_0); -- 
    maxPool4_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(21) & maxPool4_CP_346_elements(42);
      gj_maxPool4_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	70 
    -- CP-element group 41: 	74 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	82 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_update_start_
      -- CP-element group 41: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/$entry
      -- CP-element group 41: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/word_access_complete/$entry
      -- CP-element group 41: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/word_access_complete/word_0/cr
      -- 
    cr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(41), ack => ptr_deref_123_load_0_req_1); -- 
    maxPool4_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(70) & maxPool4_CP_346_elements(74) & maxPool4_CP_346_elements(78) & maxPool4_CP_346_elements(82);
      gj_maxPool4_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	16 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_sample_completed_
      -- CP-element group 42: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/word_access_start/$exit
      -- CP-element group 42: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Sample/word_access_start/word_0/ra
      -- 
    ra_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_123_load_0_ack_0, ack => maxPool4_CP_346_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	68 
    -- CP-element group 43: 	72 
    -- CP-element group 43: 	76 
    -- CP-element group 43: 	80 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_update_completed_
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/$exit
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/word_access_complete/$exit
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/ptr_deref_123_Merge/$entry
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/ptr_deref_123_Merge/$exit
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/ptr_deref_123_Merge/merge_req
      -- CP-element group 43: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_123_Update/ptr_deref_123_Merge/merge_ack
      -- 
    ca_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_123_load_0_ack_1, ack => maxPool4_CP_346_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	28 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_sample_start_
      -- CP-element group 44: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/$entry
      -- CP-element group 44: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/word_access_start/$entry
      -- CP-element group 44: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/word_access_start/word_0/rr
      -- 
    rr_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(44), ack => ptr_deref_127_load_0_req_0); -- 
    maxPool4_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(28) & maxPool4_CP_346_elements(46);
      gj_maxPool4_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	86 
    -- CP-element group 45: 	90 
    -- CP-element group 45: 	94 
    -- CP-element group 45: 	98 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_update_start_
      -- CP-element group 45: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/$entry
      -- CP-element group 45: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/word_access_complete/$entry
      -- CP-element group 45: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/word_access_complete/word_0/cr
      -- 
    cr_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(45), ack => ptr_deref_127_load_0_req_1); -- 
    maxPool4_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(86) & maxPool4_CP_346_elements(90) & maxPool4_CP_346_elements(94) & maxPool4_CP_346_elements(98);
      gj_maxPool4_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_sample_completed_
      -- CP-element group 46: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Sample/word_access_start/word_0/ra
      -- 
    ra_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_127_load_0_ack_0, ack => maxPool4_CP_346_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	84 
    -- CP-element group 47: 	88 
    -- CP-element group 47: 	92 
    -- CP-element group 47: 	96 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_update_completed_
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/$exit
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/ptr_deref_127_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/ptr_deref_127_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/ptr_deref_127_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_127_Update/ptr_deref_127_Merge/merge_ack
      -- 
    ca_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_127_load_0_ack_1, ack => maxPool4_CP_346_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_sample_start_
      -- CP-element group 48: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/word_access_start/$entry
      -- CP-element group 48: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/word_access_start/word_0/rr
      -- 
    rr_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(48), ack => ptr_deref_131_load_0_req_0); -- 
    maxPool4_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(35) & maxPool4_CP_346_elements(50);
      gj_maxPool4_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	102 
    -- CP-element group 49: 	106 
    -- CP-element group 49: 	110 
    -- CP-element group 49: 	114 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_update_start_
      -- CP-element group 49: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/$entry
      -- CP-element group 49: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/word_access_complete/$entry
      -- CP-element group 49: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/word_access_complete/word_0/$entry
      -- CP-element group 49: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/word_access_complete/word_0/cr
      -- 
    cr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(49), ack => ptr_deref_131_load_0_req_1); -- 
    maxPool4_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(102) & maxPool4_CP_346_elements(106) & maxPool4_CP_346_elements(110) & maxPool4_CP_346_elements(114);
      gj_maxPool4_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	30 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_sample_completed_
      -- CP-element group 50: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/word_access_start/$exit
      -- CP-element group 50: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Sample/word_access_start/word_0/ra
      -- 
    ra_731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_131_load_0_ack_0, ack => maxPool4_CP_346_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: 	104 
    -- CP-element group 51: 	108 
    -- CP-element group 51: 	112 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_update_completed_
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/$exit
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/word_access_complete/$exit
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/ptr_deref_131_Merge/$entry
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/ptr_deref_131_Merge/$exit
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/ptr_deref_131_Merge/merge_req
      -- CP-element group 51: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_131_Update/ptr_deref_131_Merge/merge_ack
      -- 
    ca_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_131_load_0_ack_1, ack => maxPool4_CP_346_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	39 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_95_to_assign_stmt_386/slice_136_sample_start_
      -- CP-element group 52: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Sample/rr
      -- 
    rr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(52), ack => slice_136_inst_req_0); -- 
    maxPool4_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(54);
      gj_maxPool4_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	129 
    -- CP-element group 53: 	137 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_95_to_assign_stmt_386/slice_136_update_start_
      -- CP-element group 53: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Update/$entry
      -- CP-element group 53: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Update/cr
      -- 
    cr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(53), ack => slice_136_inst_req_1); -- 
    maxPool4_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(55) & maxPool4_CP_346_elements(129) & maxPool4_CP_346_elements(137);
      gj_maxPool4_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_95_to_assign_stmt_386/slice_136_sample_completed_
      -- CP-element group 54: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Sample/ra
      -- 
    ra_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_136_inst_ack_0, ack => maxPool4_CP_346_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	127 
    -- CP-element group 55: 	135 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_95_to_assign_stmt_386/slice_136_update_completed_
      -- CP-element group 55: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Update/$exit
      -- CP-element group 55: 	 assign_stmt_95_to_assign_stmt_386/slice_136_Update/ca
      -- 
    ca_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_136_inst_ack_1, ack => maxPool4_CP_346_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_95_to_assign_stmt_386/slice_140_sample_start_
      -- CP-element group 56: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Sample/rr
      -- 
    rr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(56), ack => slice_140_inst_req_0); -- 
    maxPool4_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(58);
      gj_maxPool4_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	129 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_95_to_assign_stmt_386/slice_140_update_start_
      -- CP-element group 57: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Update/$entry
      -- CP-element group 57: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Update/cr
      -- 
    cr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(57), ack => slice_140_inst_req_1); -- 
    maxPool4_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(59) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_95_to_assign_stmt_386/slice_140_sample_completed_
      -- CP-element group 58: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Sample/$exit
      -- CP-element group 58: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Sample/ra
      -- 
    ra_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_140_inst_ack_0, ack => maxPool4_CP_346_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	127 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_95_to_assign_stmt_386/slice_140_update_completed_
      -- CP-element group 59: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Update/$exit
      -- CP-element group 59: 	 assign_stmt_95_to_assign_stmt_386/slice_140_Update/ca
      -- 
    ca_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_140_inst_ack_1, ack => maxPool4_CP_346_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_95_to_assign_stmt_386/slice_144_sample_start_
      -- CP-element group 60: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Sample/$entry
      -- CP-element group 60: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Sample/rr
      -- 
    rr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(60), ack => slice_144_inst_req_0); -- 
    maxPool4_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(62);
      gj_maxPool4_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	129 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_95_to_assign_stmt_386/slice_144_update_start_
      -- CP-element group 61: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Update/$entry
      -- CP-element group 61: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Update/cr
      -- 
    cr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(61), ack => slice_144_inst_req_1); -- 
    maxPool4_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(63) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_95_to_assign_stmt_386/slice_144_sample_completed_
      -- CP-element group 62: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Sample/ra
      -- 
    ra_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_144_inst_ack_0, ack => maxPool4_CP_346_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	127 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_95_to_assign_stmt_386/slice_144_update_completed_
      -- CP-element group 63: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Update/$exit
      -- CP-element group 63: 	 assign_stmt_95_to_assign_stmt_386/slice_144_Update/ca
      -- 
    ca_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_144_inst_ack_1, ack => maxPool4_CP_346_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_95_to_assign_stmt_386/slice_148_sample_start_
      -- CP-element group 64: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Sample/rr
      -- 
    rr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(64), ack => slice_148_inst_req_0); -- 
    maxPool4_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(66);
      gj_maxPool4_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	129 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_95_to_assign_stmt_386/slice_148_update_start_
      -- CP-element group 65: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Update/$entry
      -- CP-element group 65: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Update/cr
      -- 
    cr_802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(65), ack => slice_148_inst_req_1); -- 
    maxPool4_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(67) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_95_to_assign_stmt_386/slice_148_sample_completed_
      -- CP-element group 66: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Sample/ra
      -- 
    ra_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_148_inst_ack_0, ack => maxPool4_CP_346_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	127 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_95_to_assign_stmt_386/slice_148_update_completed_
      -- CP-element group 67: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Update/$exit
      -- CP-element group 67: 	 assign_stmt_95_to_assign_stmt_386/slice_148_Update/ca
      -- 
    ca_803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_148_inst_ack_1, ack => maxPool4_CP_346_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	43 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_95_to_assign_stmt_386/slice_152_sample_start_
      -- CP-element group 68: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Sample/$entry
      -- CP-element group 68: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Sample/rr
      -- 
    rr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(68), ack => slice_152_inst_req_0); -- 
    maxPool4_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(70);
      gj_maxPool4_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: 	129 
    -- CP-element group 69: 	137 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_95_to_assign_stmt_386/slice_152_update_start_
      -- CP-element group 69: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Update/$entry
      -- CP-element group 69: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Update/cr
      -- 
    cr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(69), ack => slice_152_inst_req_1); -- 
    maxPool4_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(71) & maxPool4_CP_346_elements(129) & maxPool4_CP_346_elements(137);
      gj_maxPool4_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	41 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_95_to_assign_stmt_386/slice_152_sample_completed_
      -- CP-element group 70: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Sample/$exit
      -- CP-element group 70: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Sample/ra
      -- 
    ra_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_152_inst_ack_0, ack => maxPool4_CP_346_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	127 
    -- CP-element group 71: 	135 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_95_to_assign_stmt_386/slice_152_update_completed_
      -- CP-element group 71: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Update/$exit
      -- CP-element group 71: 	 assign_stmt_95_to_assign_stmt_386/slice_152_Update/ca
      -- 
    ca_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_152_inst_ack_1, ack => maxPool4_CP_346_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	43 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 assign_stmt_95_to_assign_stmt_386/slice_156_sample_start_
      -- CP-element group 72: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Sample/rr
      -- 
    rr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(72), ack => slice_156_inst_req_0); -- 
    maxPool4_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(74);
      gj_maxPool4_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	129 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_95_to_assign_stmt_386/slice_156_update_start_
      -- CP-element group 73: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Update/$entry
      -- CP-element group 73: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Update/cr
      -- 
    cr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(73), ack => slice_156_inst_req_1); -- 
    maxPool4_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(75) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	41 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_95_to_assign_stmt_386/slice_156_sample_completed_
      -- CP-element group 74: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Sample/ra
      -- 
    ra_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_156_inst_ack_0, ack => maxPool4_CP_346_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	127 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_95_to_assign_stmt_386/slice_156_update_completed_
      -- CP-element group 75: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Update/$exit
      -- CP-element group 75: 	 assign_stmt_95_to_assign_stmt_386/slice_156_Update/ca
      -- 
    ca_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_156_inst_ack_1, ack => maxPool4_CP_346_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	43 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 assign_stmt_95_to_assign_stmt_386/slice_160_sample_start_
      -- CP-element group 76: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Sample/$entry
      -- CP-element group 76: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Sample/rr
      -- 
    rr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(76), ack => slice_160_inst_req_0); -- 
    maxPool4_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(78);
      gj_maxPool4_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	129 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_95_to_assign_stmt_386/slice_160_update_start_
      -- CP-element group 77: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Update/$entry
      -- CP-element group 77: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Update/cr
      -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(77), ack => slice_160_inst_req_1); -- 
    maxPool4_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(79) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_95_to_assign_stmt_386/slice_160_sample_completed_
      -- CP-element group 78: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Sample/$exit
      -- CP-element group 78: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Sample/ra
      -- 
    ra_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_160_inst_ack_0, ack => maxPool4_CP_346_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	127 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_95_to_assign_stmt_386/slice_160_update_completed_
      -- CP-element group 79: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Update/$exit
      -- CP-element group 79: 	 assign_stmt_95_to_assign_stmt_386/slice_160_Update/ca
      -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_160_inst_ack_1, ack => maxPool4_CP_346_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_95_to_assign_stmt_386/slice_164_sample_start_
      -- CP-element group 80: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Sample/$entry
      -- CP-element group 80: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Sample/rr
      -- 
    rr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(80), ack => slice_164_inst_req_0); -- 
    maxPool4_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(82);
      gj_maxPool4_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	129 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 assign_stmt_95_to_assign_stmt_386/slice_164_update_start_
      -- CP-element group 81: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Update/$entry
      -- CP-element group 81: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Update/cr
      -- 
    cr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(81), ack => slice_164_inst_req_1); -- 
    maxPool4_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(83) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	41 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_95_to_assign_stmt_386/slice_164_sample_completed_
      -- CP-element group 82: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Sample/ra
      -- 
    ra_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_164_inst_ack_0, ack => maxPool4_CP_346_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	127 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_95_to_assign_stmt_386/slice_164_update_completed_
      -- CP-element group 83: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Update/$exit
      -- CP-element group 83: 	 assign_stmt_95_to_assign_stmt_386/slice_164_Update/ca
      -- 
    ca_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_164_inst_ack_1, ack => maxPool4_CP_346_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	47 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_95_to_assign_stmt_386/slice_168_sample_start_
      -- CP-element group 84: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Sample/$entry
      -- CP-element group 84: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Sample/rr
      -- 
    rr_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(84), ack => slice_168_inst_req_0); -- 
    maxPool4_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(86);
      gj_maxPool4_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: 	129 
    -- CP-element group 85: 	137 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 assign_stmt_95_to_assign_stmt_386/slice_168_update_start_
      -- CP-element group 85: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Update/$entry
      -- CP-element group 85: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Update/cr
      -- 
    cr_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(85), ack => slice_168_inst_req_1); -- 
    maxPool4_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(87) & maxPool4_CP_346_elements(129) & maxPool4_CP_346_elements(137);
      gj_maxPool4_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	45 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_95_to_assign_stmt_386/slice_168_sample_completed_
      -- CP-element group 86: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Sample/ra
      -- 
    ra_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_168_inst_ack_0, ack => maxPool4_CP_346_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	127 
    -- CP-element group 87: 	135 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_95_to_assign_stmt_386/slice_168_update_completed_
      -- CP-element group 87: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Update/$exit
      -- CP-element group 87: 	 assign_stmt_95_to_assign_stmt_386/slice_168_Update/ca
      -- 
    ca_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_168_inst_ack_1, ack => maxPool4_CP_346_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	47 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_95_to_assign_stmt_386/slice_172_sample_start_
      -- CP-element group 88: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Sample/rr
      -- 
    rr_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(88), ack => slice_172_inst_req_0); -- 
    maxPool4_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(90);
      gj_maxPool4_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	129 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_95_to_assign_stmt_386/slice_172_update_start_
      -- CP-element group 89: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Update/$entry
      -- CP-element group 89: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Update/cr
      -- 
    cr_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(89), ack => slice_172_inst_req_1); -- 
    maxPool4_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(91) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	45 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 assign_stmt_95_to_assign_stmt_386/slice_172_sample_completed_
      -- CP-element group 90: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Sample/$exit
      -- CP-element group 90: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Sample/ra
      -- 
    ra_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_172_inst_ack_0, ack => maxPool4_CP_346_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	127 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_95_to_assign_stmt_386/slice_172_update_completed_
      -- CP-element group 91: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Update/$exit
      -- CP-element group 91: 	 assign_stmt_95_to_assign_stmt_386/slice_172_Update/ca
      -- 
    ca_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_172_inst_ack_1, ack => maxPool4_CP_346_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	47 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_95_to_assign_stmt_386/slice_176_sample_start_
      -- CP-element group 92: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Sample/rr
      -- 
    rr_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(92), ack => slice_176_inst_req_0); -- 
    maxPool4_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(94);
      gj_maxPool4_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	129 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_95_to_assign_stmt_386/slice_176_update_start_
      -- CP-element group 93: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Update/$entry
      -- CP-element group 93: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Update/cr
      -- 
    cr_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(93), ack => slice_176_inst_req_1); -- 
    maxPool4_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(95) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	45 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_95_to_assign_stmt_386/slice_176_sample_completed_
      -- CP-element group 94: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Sample/ra
      -- 
    ra_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_176_inst_ack_0, ack => maxPool4_CP_346_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	127 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_95_to_assign_stmt_386/slice_176_update_completed_
      -- CP-element group 95: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Update/$exit
      -- CP-element group 95: 	 assign_stmt_95_to_assign_stmt_386/slice_176_Update/ca
      -- 
    ca_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_176_inst_ack_1, ack => maxPool4_CP_346_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	47 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_95_to_assign_stmt_386/slice_180_sample_start_
      -- CP-element group 96: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Sample/$entry
      -- CP-element group 96: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Sample/rr
      -- 
    rr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(96), ack => slice_180_inst_req_0); -- 
    maxPool4_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(98);
      gj_maxPool4_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	129 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_95_to_assign_stmt_386/slice_180_update_start_
      -- CP-element group 97: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Update/$entry
      -- CP-element group 97: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Update/cr
      -- 
    cr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(97), ack => slice_180_inst_req_1); -- 
    maxPool4_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(99) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	45 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_95_to_assign_stmt_386/slice_180_sample_completed_
      -- CP-element group 98: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Sample/ra
      -- 
    ra_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_180_inst_ack_0, ack => maxPool4_CP_346_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	127 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 assign_stmt_95_to_assign_stmt_386/slice_180_update_completed_
      -- CP-element group 99: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Update/$exit
      -- CP-element group 99: 	 assign_stmt_95_to_assign_stmt_386/slice_180_Update/ca
      -- 
    ca_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_180_inst_ack_1, ack => maxPool4_CP_346_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	51 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_95_to_assign_stmt_386/slice_184_sample_start_
      -- CP-element group 100: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Sample/$entry
      -- CP-element group 100: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Sample/rr
      -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(100), ack => slice_184_inst_req_0); -- 
    maxPool4_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(102);
      gj_maxPool4_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	129 
    -- CP-element group 101: 	137 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 assign_stmt_95_to_assign_stmt_386/slice_184_update_start_
      -- CP-element group 101: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Update/$entry
      -- CP-element group 101: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Update/cr
      -- 
    cr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(101), ack => slice_184_inst_req_1); -- 
    maxPool4_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(103) & maxPool4_CP_346_elements(129) & maxPool4_CP_346_elements(137);
      gj_maxPool4_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 assign_stmt_95_to_assign_stmt_386/slice_184_sample_completed_
      -- CP-element group 102: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Sample/ra
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_184_inst_ack_0, ack => maxPool4_CP_346_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	127 
    -- CP-element group 103: 	135 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 assign_stmt_95_to_assign_stmt_386/slice_184_update_completed_
      -- CP-element group 103: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Update/$exit
      -- CP-element group 103: 	 assign_stmt_95_to_assign_stmt_386/slice_184_Update/ca
      -- 
    ca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_184_inst_ack_1, ack => maxPool4_CP_346_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	51 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_95_to_assign_stmt_386/slice_188_sample_start_
      -- CP-element group 104: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Sample/$entry
      -- CP-element group 104: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Sample/rr
      -- 
    rr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(104), ack => slice_188_inst_req_0); -- 
    maxPool4_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(106);
      gj_maxPool4_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	129 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_95_to_assign_stmt_386/slice_188_update_start_
      -- CP-element group 105: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Update/$entry
      -- CP-element group 105: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Update/cr
      -- 
    cr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(105), ack => slice_188_inst_req_1); -- 
    maxPool4_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(107) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	49 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_95_to_assign_stmt_386/slice_188_sample_completed_
      -- CP-element group 106: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Sample/$exit
      -- CP-element group 106: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Sample/ra
      -- 
    ra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_188_inst_ack_0, ack => maxPool4_CP_346_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	127 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_95_to_assign_stmt_386/slice_188_update_completed_
      -- CP-element group 107: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Update/$exit
      -- CP-element group 107: 	 assign_stmt_95_to_assign_stmt_386/slice_188_Update/ca
      -- 
    ca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_188_inst_ack_1, ack => maxPool4_CP_346_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	51 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 assign_stmt_95_to_assign_stmt_386/slice_192_sample_start_
      -- CP-element group 108: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Sample/rr
      -- 
    rr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(108), ack => slice_192_inst_req_0); -- 
    maxPool4_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(110);
      gj_maxPool4_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	129 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 assign_stmt_95_to_assign_stmt_386/slice_192_update_start_
      -- CP-element group 109: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Update/$entry
      -- CP-element group 109: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Update/cr
      -- 
    cr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(109), ack => slice_192_inst_req_1); -- 
    maxPool4_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(111) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 assign_stmt_95_to_assign_stmt_386/slice_192_sample_completed_
      -- CP-element group 110: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Sample/$exit
      -- CP-element group 110: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Sample/ra
      -- 
    ra_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_192_inst_ack_0, ack => maxPool4_CP_346_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	127 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 assign_stmt_95_to_assign_stmt_386/slice_192_update_completed_
      -- CP-element group 111: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Update/$exit
      -- CP-element group 111: 	 assign_stmt_95_to_assign_stmt_386/slice_192_Update/ca
      -- 
    ca_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_192_inst_ack_1, ack => maxPool4_CP_346_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	51 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 assign_stmt_95_to_assign_stmt_386/slice_196_sample_start_
      -- CP-element group 112: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Sample/$entry
      -- CP-element group 112: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Sample/rr
      -- 
    rr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(112), ack => slice_196_inst_req_0); -- 
    maxPool4_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(114);
      gj_maxPool4_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	129 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_95_to_assign_stmt_386/slice_196_update_start_
      -- CP-element group 113: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Update/$entry
      -- CP-element group 113: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Update/cr
      -- 
    cr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(113), ack => slice_196_inst_req_1); -- 
    maxPool4_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(115) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	49 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_95_to_assign_stmt_386/slice_196_sample_completed_
      -- CP-element group 114: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Sample/$exit
      -- CP-element group 114: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Sample/ra
      -- 
    ra_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_196_inst_ack_0, ack => maxPool4_CP_346_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	127 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_95_to_assign_stmt_386/slice_196_update_completed_
      -- CP-element group 115: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Update/$exit
      -- CP-element group 115: 	 assign_stmt_95_to_assign_stmt_386/slice_196_Update/ca
      -- 
    ca_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_196_inst_ack_1, ack => maxPool4_CP_346_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	120 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	121 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	121 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_request/req
      -- CP-element group 116: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_request/$entry
      -- CP-element group 116: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_sample_start_
      -- 
    req_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(116), ack => addr_of_364_final_reg_req_0); -- 
    maxPool4_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(120) & maxPool4_CP_346_elements(121);
      gj_maxPool4_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	1 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	122 
    -- CP-element group 117: 	125 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	122 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_complete/$entry
      -- CP-element group 117: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_complete/req
      -- CP-element group 117: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_update_start_
      -- 
    req_1016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(117), ack => addr_of_364_final_reg_req_1); -- 
    maxPool4_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(122) & maxPool4_CP_346_elements(125);
      gj_maxPool4_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	1 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: 	121 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_update_start
      -- CP-element group 118: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Update/$entry
      -- CP-element group 118: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Update/req
      -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(118), ack => array_obj_ref_363_index_offset_req_1); -- 
    maxPool4_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(120) & maxPool4_CP_346_elements(121);
      gj_maxPool4_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	1 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	139 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	2 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_sample_complete
      -- CP-element group 119: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Sample/$exit
      -- CP-element group 119: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Sample/ack
      -- 
    ack_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_offset_ack_0, ack => maxPool4_CP_346_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	116 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (8) 
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_base_plus_offset/sum_rename_ack
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_base_plus_offset/sum_rename_req
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_base_plus_offset/$exit
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_base_plus_offset/$entry
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_root_address_calculated
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_offset_calculated
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Update/$exit
      -- CP-element group 120: 	 assign_stmt_95_to_assign_stmt_386/array_obj_ref_363_final_index_sum_regn_Update/ack
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_offset_ack_1, ack => maxPool4_CP_346_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	116 
    -- CP-element group 121: successors 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	116 
    -- CP-element group 121: 	118 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_request/$exit
      -- CP-element group 121: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_request/ack
      -- CP-element group 121: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_sample_completed_
      -- 
    ack_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_364_final_reg_ack_0, ack => maxPool4_CP_346_elements(121)); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	117 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	117 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_complete/$exit
      -- CP-element group 122: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_complete/ack
      -- CP-element group 122: 	 assign_stmt_95_to_assign_stmt_386/addr_of_364_update_completed_
      -- 
    ack_1017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_364_final_reg_ack_1, ack => maxPool4_CP_346_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Sample/req
      -- CP-element group 123: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Sample/$entry
      -- CP-element group 123: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_sample_start_
      -- 
    req_1025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(123), ack => W_myptr5_366_delayed_8_0_366_inst_req_0); -- 
    maxPool4_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(122) & maxPool4_CP_346_elements(125);
      gj_maxPool4_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: 	133 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Update/$entry
      -- CP-element group 124: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_update_start_
      -- CP-element group 124: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Update/req
      -- 
    req_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(124), ack => W_myptr5_366_delayed_8_0_366_inst_req_1); -- 
    maxPool4_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(126) & maxPool4_CP_346_elements(133);
      gj_maxPool4_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	117 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Sample/ack
      -- CP-element group 125: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Sample/$exit
      -- CP-element group 125: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_sample_completed_
      -- 
    ack_1026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_366_delayed_8_0_366_inst_ack_0, ack => maxPool4_CP_346_elements(125)); -- 
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	131 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (19) 
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_word_addrgen/$exit
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Update/$exit
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_root_address_calculated
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_word_address_calculated
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_word_addrgen/root_register_ack
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_word_addrgen/root_register_req
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_word_addrgen/$entry
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_address_calculated
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_update_completed_
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_plus_offset/$exit
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_plus_offset/$entry
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_addr_resize/base_resize_ack
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_addr_resize/base_resize_req
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_addr_resize/$exit
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_addr_resize/$entry
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/assign_stmt_368_Update/ack
      -- CP-element group 126: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_base_address_resized
      -- 
    ack_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_366_delayed_8_0_366_inst_ack_1, ack => maxPool4_CP_346_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	55 
    -- CP-element group 127: 	59 
    -- CP-element group 127: 	63 
    -- CP-element group 127: 	67 
    -- CP-element group 127: 	71 
    -- CP-element group 127: 	75 
    -- CP-element group 127: 	79 
    -- CP-element group 127: 	83 
    -- CP-element group 127: 	87 
    -- CP-element group 127: 	91 
    -- CP-element group 127: 	95 
    -- CP-element group 127: 	99 
    -- CP-element group 127: 	103 
    -- CP-element group 127: 	107 
    -- CP-element group 127: 	111 
    -- CP-element group 127: 	115 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Sample/$entry
      -- CP-element group 127: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Sample/rr
      -- CP-element group 127: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_sample_start_
      -- 
    rr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(127), ack => CONCAT_u32_u64_381_inst_req_0); -- 
    maxPool4_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(55) & maxPool4_CP_346_elements(59) & maxPool4_CP_346_elements(63) & maxPool4_CP_346_elements(67) & maxPool4_CP_346_elements(71) & maxPool4_CP_346_elements(75) & maxPool4_CP_346_elements(79) & maxPool4_CP_346_elements(83) & maxPool4_CP_346_elements(87) & maxPool4_CP_346_elements(91) & maxPool4_CP_346_elements(95) & maxPool4_CP_346_elements(99) & maxPool4_CP_346_elements(103) & maxPool4_CP_346_elements(107) & maxPool4_CP_346_elements(111) & maxPool4_CP_346_elements(115) & maxPool4_CP_346_elements(129);
      gj_maxPool4_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Update/cr
      -- CP-element group 128: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Update/$entry
      -- CP-element group 128: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_update_start_
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(128), ack => CONCAT_u32_u64_381_inst_req_1); -- 
    maxPool4_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(130) & maxPool4_CP_346_elements(133);
      gj_maxPool4_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	53 
    -- CP-element group 129: 	57 
    -- CP-element group 129: 	61 
    -- CP-element group 129: 	65 
    -- CP-element group 129: 	69 
    -- CP-element group 129: 	73 
    -- CP-element group 129: 	77 
    -- CP-element group 129: 	81 
    -- CP-element group 129: 	85 
    -- CP-element group 129: 	89 
    -- CP-element group 129: 	93 
    -- CP-element group 129: 	97 
    -- CP-element group 129: 	101 
    -- CP-element group 129: 	105 
    -- CP-element group 129: 	109 
    -- CP-element group 129: 	113 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Sample/ra
      -- CP-element group 129: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Sample/$exit
      -- CP-element group 129: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_sample_completed_
      -- 
    ra_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_381_inst_ack_0, ack => maxPool4_CP_346_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Update/ca
      -- CP-element group 130: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_Update/$exit
      -- CP-element group 130: 	 assign_stmt_95_to_assign_stmt_386/CONCAT_u32_u64_381_update_completed_
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_381_inst_ack_1, ack => maxPool4_CP_346_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	126 
    -- CP-element group 131: 	130 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (9) 
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/word_access_start/$entry
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/ptr_deref_370_Split/split_ack
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/ptr_deref_370_Split/split_req
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_sample_start_
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/ptr_deref_370_Split/$exit
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/ptr_deref_370_Split/$entry
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/$entry
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/word_access_start/word_0/rr
      -- CP-element group 131: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/word_access_start/word_0/$entry
      -- 
    rr_1083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(131), ack => ptr_deref_370_store_0_req_0); -- 
    maxPool4_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(126) & maxPool4_CP_346_elements(130) & maxPool4_CP_346_elements(133);
      gj_maxPool4_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/$entry
      -- CP-element group 132: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/word_access_complete/word_0/cr
      -- CP-element group 132: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/word_access_complete/word_0/$entry
      -- CP-element group 132: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_update_start_
      -- CP-element group 132: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/word_access_complete/$entry
      -- 
    cr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(132), ack => ptr_deref_370_store_0_req_1); -- 
    maxPool4_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(134);
      gj_maxPool4_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	124 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/word_access_start/$exit
      -- CP-element group 133: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_sample_completed_
      -- CP-element group 133: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/$exit
      -- CP-element group 133: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/word_access_start/word_0/ra
      -- CP-element group 133: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Sample/word_access_start/word_0/$exit
      -- 
    ra_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_370_store_0_ack_0, ack => maxPool4_CP_346_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	139 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/$exit
      -- CP-element group 134: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_update_completed_
      -- CP-element group 134: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/word_access_complete/word_0/ca
      -- CP-element group 134: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/word_access_complete/word_0/$exit
      -- CP-element group 134: 	 assign_stmt_95_to_assign_stmt_386/ptr_deref_370_Update/word_access_complete/$exit
      -- 
    ca_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_370_store_0_ack_1, ack => maxPool4_CP_346_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	55 
    -- CP-element group 135: 	71 
    -- CP-element group 135: 	87 
    -- CP-element group 135: 	103 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Sample/rr
      -- CP-element group 135: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Sample/$entry
      -- CP-element group 135: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_sample_start_
      -- 
    rr_1103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(135), ack => type_cast_385_inst_req_0); -- 
    maxPool4_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(55) & maxPool4_CP_346_elements(71) & maxPool4_CP_346_elements(87) & maxPool4_CP_346_elements(103) & maxPool4_CP_346_elements(137);
      gj_maxPool4_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	7 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Update/cr
      -- CP-element group 136: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_update_start_
      -- CP-element group 136: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Update/$entry
      -- 
    cr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(136), ack => type_cast_385_inst_req_1); -- 
    maxPool4_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(7) & maxPool4_CP_346_elements(138);
      gj_maxPool4_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	53 
    -- CP-element group 137: 	69 
    -- CP-element group 137: 	85 
    -- CP-element group 137: 	101 
    -- CP-element group 137: 	135 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Sample/ra
      -- CP-element group 137: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Sample/$exit
      -- CP-element group 137: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_sample_completed_
      -- 
    ra_1104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_385_inst_ack_0, ack => maxPool4_CP_346_elements(137)); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Update/ca
      -- CP-element group 138: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_update_completed_
      -- CP-element group 138: 	 assign_stmt_95_to_assign_stmt_386/type_cast_385_Update/$exit
      -- 
    ca_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_385_inst_ack_1, ack => maxPool4_CP_346_elements(138)); -- 
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	11 
    -- CP-element group 139: 	18 
    -- CP-element group 139: 	25 
    -- CP-element group 139: 	32 
    -- CP-element group 139: 	119 
    -- CP-element group 139: 	134 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	146 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 assign_stmt_95_to_assign_stmt_386/$exit
      -- 
    maxPool4_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(11) & maxPool4_CP_346_elements(18) & maxPool4_CP_346_elements(25) & maxPool4_CP_346_elements(32) & maxPool4_CP_346_elements(119) & maxPool4_CP_346_elements(134) & maxPool4_CP_346_elements(138);
      gj_maxPool4_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  place  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	2 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 addr_update_enable
      -- 
    maxPool4_CP_346_elements(140) <= maxPool4_CP_346_elements(2);
    -- CP-element group 141:  place  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	3 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 addr1_update_enable
      -- 
    maxPool4_CP_346_elements(141) <= maxPool4_CP_346_elements(3);
    -- CP-element group 142:  place  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	4 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 addr2_update_enable
      -- 
    maxPool4_CP_346_elements(142) <= maxPool4_CP_346_elements(4);
    -- CP-element group 143:  place  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	5 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 addr3_update_enable
      -- 
    maxPool4_CP_346_elements(143) <= maxPool4_CP_346_elements(5);
    -- CP-element group 144:  place  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	6 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 addr4_update_enable
      -- 
    maxPool4_CP_346_elements(144) <= maxPool4_CP_346_elements(6);
    -- CP-element group 145:  place  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	7 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 output_update_enable
      -- 
    -- CP-element group 146:  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	139 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 $exit
      -- 
    maxPool4_CP_346_elements(146) <= maxPool4_CP_346_elements(139);
    --  hookup: inputs to control-path 
    maxPool4_CP_346_elements(145) <= output_update_enable;
    -- hookup: output from control-path 
    addr4_update_enable <= maxPool4_CP_346_elements(144);
    addr_update_enable <= maxPool4_CP_346_elements(140);
    addr3_update_enable <= maxPool4_CP_346_elements(143);
    addr2_update_enable <= maxPool4_CP_346_elements(142);
    addr1_update_enable <= maxPool4_CP_346_elements(141);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_375_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_380_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_381_wire : std_logic_vector(63 downto 0);
    signal R_addr1_92_resized : std_logic_vector(13 downto 0);
    signal R_addr1_92_scaled : std_logic_vector(13 downto 0);
    signal R_addr2_99_resized : std_logic_vector(13 downto 0);
    signal R_addr2_99_scaled : std_logic_vector(13 downto 0);
    signal R_addr3_106_resized : std_logic_vector(13 downto 0);
    signal R_addr3_106_scaled : std_logic_vector(13 downto 0);
    signal R_addr4_113_resized : std_logic_vector(13 downto 0);
    signal R_addr4_113_scaled : std_logic_vector(13 downto 0);
    signal R_addr_362_resized : std_logic_vector(13 downto 0);
    signal R_addr_362_scaled : std_logic_vector(13 downto 0);
    signal SGT_i16_u1_266_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_274_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_282_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_290_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_298_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_306_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_314_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_322_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_330_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_338_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_346_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_354_wire : std_logic_vector(0 downto 0);
    signal a11_202 : std_logic_vector(15 downto 0);
    signal a12_206 : std_logic_vector(15 downto 0);
    signal a13_210 : std_logic_vector(15 downto 0);
    signal a14_214 : std_logic_vector(15 downto 0);
    signal a21_218 : std_logic_vector(15 downto 0);
    signal a22_222 : std_logic_vector(15 downto 0);
    signal a23_226 : std_logic_vector(15 downto 0);
    signal a24_230 : std_logic_vector(15 downto 0);
    signal a31_234 : std_logic_vector(15 downto 0);
    signal a32_238 : std_logic_vector(15 downto 0);
    signal a33_242 : std_logic_vector(15 downto 0);
    signal a34_246 : std_logic_vector(15 downto 0);
    signal a41_250 : std_logic_vector(15 downto 0);
    signal a42_254 : std_logic_vector(15 downto 0);
    signal a43_258 : std_logic_vector(15 downto 0);
    signal a44_262 : std_logic_vector(15 downto 0);
    signal array_obj_ref_100_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_100_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_100_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_100_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_100_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_100_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_107_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_107_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_107_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_107_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_107_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_107_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_114_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_114_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_114_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_114_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_114_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_114_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_root_address : std_logic_vector(13 downto 0);
    signal c1_120 : std_logic_vector(63 downto 0);
    signal c2_124 : std_logic_vector(63 downto 0);
    signal c3_128 : std_logic_vector(63 downto 0);
    signal c4_132 : std_logic_vector(63 downto 0);
    signal myptr1_95 : std_logic_vector(31 downto 0);
    signal myptr2_102 : std_logic_vector(31 downto 0);
    signal myptr3_109 : std_logic_vector(31 downto 0);
    signal myptr4_116 : std_logic_vector(31 downto 0);
    signal myptr5_365 : std_logic_vector(31 downto 0);
    signal myptr5_366_delayed_8_0_368 : std_logic_vector(31 downto 0);
    signal out1_286 : std_logic_vector(15 downto 0);
    signal out2_310 : std_logic_vector(15 downto 0);
    signal out3_334 : std_logic_vector(15 downto 0);
    signal out4_358 : std_logic_vector(15 downto 0);
    signal ptr_deref_119_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_119_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_119_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_119_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_119_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_123_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_123_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_123_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_123_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_123_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_127_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_127_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_127_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_127_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_127_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_131_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_131_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_131_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_131_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_131_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_370_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_370_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_370_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_370_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_370_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_370_word_offset_0 : std_logic_vector(13 downto 0);
    signal sliced_v11_137 : std_logic_vector(15 downto 0);
    signal sliced_v12_141 : std_logic_vector(15 downto 0);
    signal sliced_v13_145 : std_logic_vector(15 downto 0);
    signal sliced_v14_149 : std_logic_vector(15 downto 0);
    signal sliced_v21_153 : std_logic_vector(15 downto 0);
    signal sliced_v22_157 : std_logic_vector(15 downto 0);
    signal sliced_v23_161 : std_logic_vector(15 downto 0);
    signal sliced_v24_165 : std_logic_vector(15 downto 0);
    signal sliced_v31_169 : std_logic_vector(15 downto 0);
    signal sliced_v32_173 : std_logic_vector(15 downto 0);
    signal sliced_v33_177 : std_logic_vector(15 downto 0);
    signal sliced_v34_181 : std_logic_vector(15 downto 0);
    signal sliced_v41_185 : std_logic_vector(15 downto 0);
    signal sliced_v42_189 : std_logic_vector(15 downto 0);
    signal sliced_v43_193 : std_logic_vector(15 downto 0);
    signal sliced_v44_197 : std_logic_vector(15 downto 0);
    signal t11_270 : std_logic_vector(15 downto 0);
    signal t12_278 : std_logic_vector(15 downto 0);
    signal t21_294 : std_logic_vector(15 downto 0);
    signal t22_302 : std_logic_vector(15 downto 0);
    signal t31_318 : std_logic_vector(15 downto 0);
    signal t32_326 : std_logic_vector(15 downto 0);
    signal t41_342 : std_logic_vector(15 downto 0);
    signal t42_350 : std_logic_vector(15 downto 0);
    signal type_cast_372_wire : std_logic_vector(15 downto 0);
    signal type_cast_374_wire : std_logic_vector(15 downto 0);
    signal type_cast_377_wire : std_logic_vector(15 downto 0);
    signal type_cast_379_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_100_constant_part_of_offset <= "00000000000000";
    array_obj_ref_100_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_100_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_100_resized_base_address <= "00000000000000";
    array_obj_ref_107_constant_part_of_offset <= "00000000000000";
    array_obj_ref_107_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_107_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_107_resized_base_address <= "00000000000000";
    array_obj_ref_114_constant_part_of_offset <= "00000000000000";
    array_obj_ref_114_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_114_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_114_resized_base_address <= "00000000000000";
    array_obj_ref_363_constant_part_of_offset <= "00000000000000";
    array_obj_ref_363_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_363_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_363_resized_base_address <= "00000000000000";
    array_obj_ref_93_constant_part_of_offset <= "00000000000000";
    array_obj_ref_93_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_93_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_93_resized_base_address <= "00000000000000";
    ptr_deref_119_word_offset_0 <= "00000000000000";
    ptr_deref_123_word_offset_0 <= "00000000000000";
    ptr_deref_127_word_offset_0 <= "00000000000000";
    ptr_deref_131_word_offset_0 <= "00000000000000";
    ptr_deref_370_word_offset_0 <= "00000000000000";
    -- flow-through select operator MUX_269_inst
    t11_270 <= a11_202 when (SGT_i16_u1_266_wire(0) /=  '0') else a21_218;
    -- flow-through select operator MUX_277_inst
    t12_278 <= a31_234 when (SGT_i16_u1_274_wire(0) /=  '0') else a41_250;
    -- flow-through select operator MUX_285_inst
    out1_286 <= t11_270 when (SGT_i16_u1_282_wire(0) /=  '0') else t12_278;
    -- flow-through select operator MUX_293_inst
    t21_294 <= a12_206 when (SGT_i16_u1_290_wire(0) /=  '0') else a22_222;
    -- flow-through select operator MUX_301_inst
    t22_302 <= a32_238 when (SGT_i16_u1_298_wire(0) /=  '0') else a42_254;
    -- flow-through select operator MUX_309_inst
    out2_310 <= t21_294 when (SGT_i16_u1_306_wire(0) /=  '0') else t22_302;
    -- flow-through select operator MUX_317_inst
    t31_318 <= a13_210 when (SGT_i16_u1_314_wire(0) /=  '0') else a23_226;
    -- flow-through select operator MUX_325_inst
    t32_326 <= a33_242 when (SGT_i16_u1_322_wire(0) /=  '0') else a43_258;
    -- flow-through select operator MUX_333_inst
    out3_334 <= t31_318 when (SGT_i16_u1_330_wire(0) /=  '0') else t32_326;
    -- flow-through select operator MUX_341_inst
    t41_342 <= a14_214 when (SGT_i16_u1_338_wire(0) /=  '0') else a24_230;
    -- flow-through select operator MUX_349_inst
    t42_350 <= a34_246 when (SGT_i16_u1_346_wire(0) /=  '0') else a44_262;
    -- flow-through select operator MUX_357_inst
    out4_358 <= t41_342 when (SGT_i16_u1_354_wire(0) /=  '0') else t42_350;
    slice_136_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_136_inst_req_0;
      slice_136_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_136_inst_req_1;
      slice_136_inst_ack_1<= update_ack(0);
      slice_136_inst: SliceSplitProtocol generic map(name => "slice_136_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_120, dout => sliced_v11_137, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_140_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_140_inst_req_0;
      slice_140_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_140_inst_req_1;
      slice_140_inst_ack_1<= update_ack(0);
      slice_140_inst: SliceSplitProtocol generic map(name => "slice_140_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_120, dout => sliced_v12_141, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_144_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_144_inst_req_0;
      slice_144_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_144_inst_req_1;
      slice_144_inst_ack_1<= update_ack(0);
      slice_144_inst: SliceSplitProtocol generic map(name => "slice_144_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_120, dout => sliced_v13_145, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_148_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_148_inst_req_0;
      slice_148_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_148_inst_req_1;
      slice_148_inst_ack_1<= update_ack(0);
      slice_148_inst: SliceSplitProtocol generic map(name => "slice_148_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_120, dout => sliced_v14_149, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_152_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_152_inst_req_0;
      slice_152_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_152_inst_req_1;
      slice_152_inst_ack_1<= update_ack(0);
      slice_152_inst: SliceSplitProtocol generic map(name => "slice_152_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_124, dout => sliced_v21_153, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_156_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_156_inst_req_0;
      slice_156_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_156_inst_req_1;
      slice_156_inst_ack_1<= update_ack(0);
      slice_156_inst: SliceSplitProtocol generic map(name => "slice_156_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_124, dout => sliced_v22_157, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_160_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_160_inst_req_0;
      slice_160_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_160_inst_req_1;
      slice_160_inst_ack_1<= update_ack(0);
      slice_160_inst: SliceSplitProtocol generic map(name => "slice_160_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_124, dout => sliced_v23_161, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_164_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_164_inst_req_0;
      slice_164_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_164_inst_req_1;
      slice_164_inst_ack_1<= update_ack(0);
      slice_164_inst: SliceSplitProtocol generic map(name => "slice_164_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_124, dout => sliced_v24_165, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_168_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_168_inst_req_0;
      slice_168_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_168_inst_req_1;
      slice_168_inst_ack_1<= update_ack(0);
      slice_168_inst: SliceSplitProtocol generic map(name => "slice_168_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_128, dout => sliced_v31_169, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_172_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_172_inst_req_0;
      slice_172_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_172_inst_req_1;
      slice_172_inst_ack_1<= update_ack(0);
      slice_172_inst: SliceSplitProtocol generic map(name => "slice_172_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_128, dout => sliced_v32_173, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_176_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_176_inst_req_0;
      slice_176_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_176_inst_req_1;
      slice_176_inst_ack_1<= update_ack(0);
      slice_176_inst: SliceSplitProtocol generic map(name => "slice_176_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_128, dout => sliced_v33_177, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_180_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_180_inst_req_0;
      slice_180_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_180_inst_req_1;
      slice_180_inst_ack_1<= update_ack(0);
      slice_180_inst: SliceSplitProtocol generic map(name => "slice_180_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_128, dout => sliced_v34_181, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_184_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_184_inst_req_0;
      slice_184_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_184_inst_req_1;
      slice_184_inst_ack_1<= update_ack(0);
      slice_184_inst: SliceSplitProtocol generic map(name => "slice_184_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_132, dout => sliced_v41_185, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_188_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_188_inst_req_0;
      slice_188_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_188_inst_req_1;
      slice_188_inst_ack_1<= update_ack(0);
      slice_188_inst: SliceSplitProtocol generic map(name => "slice_188_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_132, dout => sliced_v42_189, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_192_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_192_inst_req_0;
      slice_192_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_192_inst_req_1;
      slice_192_inst_ack_1<= update_ack(0);
      slice_192_inst: SliceSplitProtocol generic map(name => "slice_192_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_132, dout => sliced_v43_193, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_196_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_196_inst_req_0;
      slice_196_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_196_inst_req_1;
      slice_196_inst_ack_1<= update_ack(0);
      slice_196_inst: SliceSplitProtocol generic map(name => "slice_196_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_132, dout => sliced_v44_197, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_myptr5_366_delayed_8_0_366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr5_366_delayed_8_0_366_inst_req_0;
      W_myptr5_366_delayed_8_0_366_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr5_366_delayed_8_0_366_inst_req_1;
      W_myptr5_366_delayed_8_0_366_inst_ack_1<= rack(0);
      W_myptr5_366_delayed_8_0_366_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr5_366_delayed_8_0_366_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr5_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_366_delayed_8_0_368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_101_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_101_final_reg_req_0;
      addr_of_101_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_101_final_reg_req_1;
      addr_of_101_final_reg_ack_1<= rack(0);
      addr_of_101_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_101_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_100_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr2_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_108_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_108_final_reg_req_0;
      addr_of_108_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_108_final_reg_req_1;
      addr_of_108_final_reg_ack_1<= rack(0);
      addr_of_108_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_108_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_107_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr3_109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_115_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_115_final_reg_req_0;
      addr_of_115_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_115_final_reg_req_1;
      addr_of_115_final_reg_ack_1<= rack(0);
      addr_of_115_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_115_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_114_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr4_116,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_364_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_364_final_reg_req_0;
      addr_of_364_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_364_final_reg_req_1;
      addr_of_364_final_reg_ack_1<= rack(0);
      addr_of_364_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_364_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_363_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_94_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_94_final_reg_req_0;
      addr_of_94_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_94_final_reg_req_1;
      addr_of_94_final_reg_ack_1<= rack(0);
      addr_of_94_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_94_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_93_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr1_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_201_inst
    process(sliced_v11_137) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v11_137(15 downto 0);
      a11_202 <= tmp_var; -- 
    end process;
    -- interlock type_cast_205_inst
    process(sliced_v12_141) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v12_141(15 downto 0);
      a12_206 <= tmp_var; -- 
    end process;
    -- interlock type_cast_209_inst
    process(sliced_v13_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v13_145(15 downto 0);
      a13_210 <= tmp_var; -- 
    end process;
    -- interlock type_cast_213_inst
    process(sliced_v14_149) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v14_149(15 downto 0);
      a14_214 <= tmp_var; -- 
    end process;
    -- interlock type_cast_217_inst
    process(sliced_v21_153) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v21_153(15 downto 0);
      a21_218 <= tmp_var; -- 
    end process;
    -- interlock type_cast_221_inst
    process(sliced_v22_157) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v22_157(15 downto 0);
      a22_222 <= tmp_var; -- 
    end process;
    -- interlock type_cast_225_inst
    process(sliced_v23_161) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v23_161(15 downto 0);
      a23_226 <= tmp_var; -- 
    end process;
    -- interlock type_cast_229_inst
    process(sliced_v24_165) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v24_165(15 downto 0);
      a24_230 <= tmp_var; -- 
    end process;
    -- interlock type_cast_233_inst
    process(sliced_v31_169) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v31_169(15 downto 0);
      a31_234 <= tmp_var; -- 
    end process;
    -- interlock type_cast_237_inst
    process(sliced_v32_173) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v32_173(15 downto 0);
      a32_238 <= tmp_var; -- 
    end process;
    -- interlock type_cast_241_inst
    process(sliced_v33_177) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v33_177(15 downto 0);
      a33_242 <= tmp_var; -- 
    end process;
    -- interlock type_cast_245_inst
    process(sliced_v34_181) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v34_181(15 downto 0);
      a34_246 <= tmp_var; -- 
    end process;
    -- interlock type_cast_249_inst
    process(sliced_v41_185) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v41_185(15 downto 0);
      a41_250 <= tmp_var; -- 
    end process;
    -- interlock type_cast_253_inst
    process(sliced_v42_189) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v42_189(15 downto 0);
      a42_254 <= tmp_var; -- 
    end process;
    -- interlock type_cast_257_inst
    process(sliced_v43_193) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v43_193(15 downto 0);
      a43_258 <= tmp_var; -- 
    end process;
    -- interlock type_cast_261_inst
    process(sliced_v44_197) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v44_197(15 downto 0);
      a44_262 <= tmp_var; -- 
    end process;
    -- interlock type_cast_372_inst
    process(out1_286) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out1_286(15 downto 0);
      type_cast_372_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_374_inst
    process(out2_310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out2_310(15 downto 0);
      type_cast_374_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_377_inst
    process(out3_334) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out3_334(15 downto 0);
      type_cast_377_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_379_inst
    process(out4_358) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out4_358(15 downto 0);
      type_cast_379_wire <= tmp_var; -- 
    end process;
    type_cast_385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_385_inst_req_0;
      type_cast_385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_385_inst_req_1;
      type_cast_385_inst_ack_1<= rack(0);
      type_cast_385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out1_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_100_index_1_rename
    process(R_addr2_99_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_99_resized;
      ov(13 downto 0) := iv;
      R_addr2_99_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_100_index_1_resize
    process(addr2_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_buffer;
      ov := iv(13 downto 0);
      R_addr2_99_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_100_root_address_inst
    process(array_obj_ref_100_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_100_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_100_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_107_index_1_rename
    process(R_addr3_106_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_106_resized;
      ov(13 downto 0) := iv;
      R_addr3_106_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_107_index_1_resize
    process(addr3_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_buffer;
      ov := iv(13 downto 0);
      R_addr3_106_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_107_root_address_inst
    process(array_obj_ref_107_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_107_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_107_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_114_index_1_rename
    process(R_addr4_113_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr4_113_resized;
      ov(13 downto 0) := iv;
      R_addr4_113_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_114_index_1_resize
    process(addr4_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr4_buffer;
      ov := iv(13 downto 0);
      R_addr4_113_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_114_root_address_inst
    process(array_obj_ref_114_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_114_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_114_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_index_1_rename
    process(R_addr_362_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_362_resized;
      ov(13 downto 0) := iv;
      R_addr_362_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_362_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_root_address_inst
    process(array_obj_ref_363_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_363_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_363_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_index_1_rename
    process(R_addr1_92_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_92_resized;
      ov(13 downto 0) := iv;
      R_addr1_92_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_index_1_resize
    process(addr1_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_buffer;
      ov := iv(13 downto 0);
      R_addr1_92_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_root_address_inst
    process(array_obj_ref_93_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_93_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_93_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_119_addr_0
    process(ptr_deref_119_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_119_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_119_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_119_base_resize
    process(myptr1_95) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr1_95;
      ov := iv(13 downto 0);
      ptr_deref_119_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_119_gather_scatter
    process(ptr_deref_119_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_119_data_0;
      ov(63 downto 0) := iv;
      c1_120 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_119_root_address_inst
    process(ptr_deref_119_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_119_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_119_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_addr_0
    process(ptr_deref_123_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_123_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_123_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_base_resize
    process(myptr2_102) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr2_102;
      ov := iv(13 downto 0);
      ptr_deref_123_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_gather_scatter
    process(ptr_deref_123_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_123_data_0;
      ov(63 downto 0) := iv;
      c2_124 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_root_address_inst
    process(ptr_deref_123_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_123_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_123_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_127_addr_0
    process(ptr_deref_127_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_127_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_127_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_127_base_resize
    process(myptr3_109) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr3_109;
      ov := iv(13 downto 0);
      ptr_deref_127_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_127_gather_scatter
    process(ptr_deref_127_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_127_data_0;
      ov(63 downto 0) := iv;
      c3_128 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_127_root_address_inst
    process(ptr_deref_127_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_127_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_127_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_131_addr_0
    process(ptr_deref_131_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_131_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_131_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_131_base_resize
    process(myptr4_116) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr4_116;
      ov := iv(13 downto 0);
      ptr_deref_131_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_131_gather_scatter
    process(ptr_deref_131_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_131_data_0;
      ov(63 downto 0) := iv;
      c4_132 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_131_root_address_inst
    process(ptr_deref_131_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_131_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_131_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_addr_0
    process(ptr_deref_370_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_370_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_370_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_base_resize
    process(myptr5_366_delayed_8_0_368) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr5_366_delayed_8_0_368;
      ov := iv(13 downto 0);
      ptr_deref_370_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_gather_scatter
    process(CONCAT_u32_u64_381_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_381_wire;
      ov(63 downto 0) := iv;
      ptr_deref_370_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_root_address_inst
    process(ptr_deref_370_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_370_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_370_root_address <= ov(13 downto 0);
      --
    end process;
    -- binary operator CONCAT_u16_u32_375_inst
    process(type_cast_372_wire, type_cast_374_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_372_wire, type_cast_374_wire, tmp_var);
      CONCAT_u16_u32_375_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_380_inst
    process(type_cast_377_wire, type_cast_379_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_377_wire, type_cast_379_wire, tmp_var);
      CONCAT_u16_u32_380_wire <= tmp_var; --
    end process;
    -- shared split operator group (2) : CONCAT_u32_u64_381_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_375_wire & CONCAT_u16_u32_380_wire;
      CONCAT_u32_u64_381_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_381_inst_req_0;
      CONCAT_u32_u64_381_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_381_inst_req_1;
      CONCAT_u32_u64_381_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator SGT_i16_u1_266_inst
    process(a11_202, a21_218) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a11_202, a21_218, tmp_var);
      SGT_i16_u1_266_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_274_inst
    process(a31_234, a41_250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a31_234, a41_250, tmp_var);
      SGT_i16_u1_274_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_282_inst
    process(t11_270, t12_278) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t11_270, t12_278, tmp_var);
      SGT_i16_u1_282_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_290_inst
    process(a12_206, a22_222) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a12_206, a22_222, tmp_var);
      SGT_i16_u1_290_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_298_inst
    process(a32_238, a42_254) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a32_238, a42_254, tmp_var);
      SGT_i16_u1_298_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_306_inst
    process(t21_294, t22_302) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t21_294, t22_302, tmp_var);
      SGT_i16_u1_306_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_314_inst
    process(a13_210, a23_226) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a13_210, a23_226, tmp_var);
      SGT_i16_u1_314_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_322_inst
    process(a33_242, a43_258) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a33_242, a43_258, tmp_var);
      SGT_i16_u1_322_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_330_inst
    process(t31_318, t32_326) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t31_318, t32_326, tmp_var);
      SGT_i16_u1_330_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_338_inst
    process(a14_214, a24_230) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a14_214, a24_230, tmp_var);
      SGT_i16_u1_338_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_346_inst
    process(a34_246, a44_262) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a34_246, a44_262, tmp_var);
      SGT_i16_u1_346_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_354_inst
    process(t41_342, t42_350) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t41_342, t42_350, tmp_var);
      SGT_i16_u1_354_wire <= tmp_var; --
    end process;
    -- shared split operator group (15) : array_obj_ref_100_index_offset 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr2_99_scaled;
      array_obj_ref_100_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_100_index_offset_req_0;
      array_obj_ref_100_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_100_index_offset_req_1;
      array_obj_ref_100_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : array_obj_ref_107_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr3_106_scaled;
      array_obj_ref_107_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_107_index_offset_req_0;
      array_obj_ref_107_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_107_index_offset_req_1;
      array_obj_ref_107_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : array_obj_ref_114_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr4_113_scaled;
      array_obj_ref_114_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_114_index_offset_req_0;
      array_obj_ref_114_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_114_index_offset_req_1;
      array_obj_ref_114_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : array_obj_ref_363_index_offset 
    ApIntAdd_group_18: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_362_scaled;
      array_obj_ref_363_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_363_index_offset_req_0;
      array_obj_ref_363_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_363_index_offset_req_1;
      array_obj_ref_363_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_18_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : array_obj_ref_93_index_offset 
    ApIntAdd_group_19: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr1_92_scaled;
      array_obj_ref_93_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_93_index_offset_req_0;
      array_obj_ref_93_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_93_index_offset_req_1;
      array_obj_ref_93_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_19_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared load operator group (0) : ptr_deref_119_load_0 ptr_deref_123_load_0 ptr_deref_127_load_0 ptr_deref_131_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_119_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_123_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_127_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_131_load_0_req_0;
      ptr_deref_119_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_123_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_127_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_131_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_119_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_123_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_127_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_131_load_0_req_1;
      ptr_deref_119_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_123_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_127_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_131_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_119_word_address_0 & ptr_deref_123_word_address_0 & ptr_deref_127_word_address_0 & ptr_deref_131_word_address_0;
      ptr_deref_119_data_0 <= data_out(255 downto 192);
      ptr_deref_123_data_0 <= data_out(191 downto 128);
      ptr_deref_127_data_0 <= data_out(127 downto 64);
      ptr_deref_131_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_370_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_370_store_0_req_0;
      ptr_deref_370_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_370_store_0_req_1;
      ptr_deref_370_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_370_word_address_0;
      data_in <= ptr_deref_370_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end maxPool4_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_1116_start: Boolean;
  signal sendB_CP_1116_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_504_inst_req_0 : boolean;
  signal addr_of_454_final_reg_req_0 : boolean;
  signal addr_of_454_final_reg_ack_0 : boolean;
  signal ptr_deref_458_load_0_req_1 : boolean;
  signal ptr_deref_458_load_0_ack_1 : boolean;
  signal type_cast_424_inst_req_1 : boolean;
  signal type_cast_424_inst_ack_1 : boolean;
  signal type_cast_511_inst_req_0 : boolean;
  signal addr_of_454_final_reg_req_1 : boolean;
  signal addr_of_454_final_reg_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_506_inst_req_1 : boolean;
  signal type_cast_424_inst_req_0 : boolean;
  signal type_cast_511_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_506_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_506_inst_ack_0 : boolean;
  signal if_stmt_397_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_506_inst_ack_1 : boolean;
  signal type_cast_424_inst_ack_0 : boolean;
  signal type_cast_511_inst_req_1 : boolean;
  signal type_cast_504_inst_ack_0 : boolean;
  signal array_obj_ref_453_index_offset_req_1 : boolean;
  signal if_stmt_397_branch_ack_1 : boolean;
  signal if_stmt_397_branch_ack_0 : boolean;
  signal ptr_deref_458_load_0_req_0 : boolean;
  signal array_obj_ref_453_index_offset_ack_1 : boolean;
  signal array_obj_ref_453_index_offset_req_0 : boolean;
  signal ptr_deref_458_load_0_ack_0 : boolean;
  signal array_obj_ref_453_index_offset_ack_0 : boolean;
  signal type_cast_504_inst_req_1 : boolean;
  signal type_cast_504_inst_ack_1 : boolean;
  signal type_cast_511_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_513_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_513_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_513_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_513_inst_ack_1 : boolean;
  signal type_cast_518_inst_req_0 : boolean;
  signal type_cast_518_inst_ack_0 : boolean;
  signal type_cast_518_inst_req_1 : boolean;
  signal type_cast_518_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_520_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_520_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_520_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_520_inst_ack_1 : boolean;
  signal type_cast_525_inst_req_0 : boolean;
  signal type_cast_525_inst_ack_0 : boolean;
  signal type_cast_525_inst_req_1 : boolean;
  signal type_cast_525_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_527_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_527_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_527_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_527_inst_ack_1 : boolean;
  signal type_cast_532_inst_req_0 : boolean;
  signal type_cast_532_inst_ack_0 : boolean;
  signal type_cast_532_inst_req_1 : boolean;
  signal type_cast_532_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_534_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_534_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_534_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_534_inst_ack_1 : boolean;
  signal type_cast_539_inst_req_0 : boolean;
  signal type_cast_539_inst_ack_0 : boolean;
  signal type_cast_539_inst_req_1 : boolean;
  signal type_cast_539_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_ack_1 : boolean;
  signal type_cast_546_inst_req_0 : boolean;
  signal type_cast_546_inst_ack_0 : boolean;
  signal type_cast_546_inst_req_1 : boolean;
  signal type_cast_546_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_548_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_548_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_548_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_548_inst_ack_1 : boolean;
  signal type_cast_553_inst_req_0 : boolean;
  signal type_cast_553_inst_ack_0 : boolean;
  signal type_cast_553_inst_req_1 : boolean;
  signal type_cast_553_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_555_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_555_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_555_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_555_inst_ack_1 : boolean;
  signal if_stmt_569_branch_req_0 : boolean;
  signal if_stmt_569_branch_ack_1 : boolean;
  signal if_stmt_569_branch_ack_0 : boolean;
  signal phi_stmt_441_req_0 : boolean;
  signal type_cast_447_inst_req_0 : boolean;
  signal type_cast_447_inst_ack_0 : boolean;
  signal type_cast_447_inst_req_1 : boolean;
  signal type_cast_447_inst_ack_1 : boolean;
  signal phi_stmt_441_req_1 : boolean;
  signal phi_stmt_441_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_1116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_1116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_1116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_1116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_1116: Block -- control-path 
    signal sendB_CP_1116_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendB_CP_1116_elements(0) <= sendB_CP_1116_start;
    sendB_CP_1116_symbol <= sendB_CP_1116_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_390/assign_stmt_396/$entry
      -- CP-element group 0: 	 branch_block_stmt_390/assign_stmt_396/$exit
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_390/R_cmp76_398_place
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397_else_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_390/$entry
      -- CP-element group 0: 	 branch_block_stmt_390/branch_block_stmt_390__entry__
      -- CP-element group 0: 	 branch_block_stmt_390/assign_stmt_396__entry__
      -- CP-element group 0: 	 branch_block_stmt_390/assign_stmt_396__exit__
      -- CP-element group 0: 	 branch_block_stmt_390/if_stmt_397__entry__
      -- 
    branch_req_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(0), ack => if_stmt_397_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_390/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_390/if_stmt_397_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_390/if_stmt_397_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/$entry
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_update_start_
      -- CP-element group 1: 	 branch_block_stmt_390/merge_stmt_403__exit__
      -- CP-element group 1: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438__entry__
      -- CP-element group 1: 	 branch_block_stmt_390/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_390/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_390/merge_stmt_403_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_390/merge_stmt_403_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_390/merge_stmt_403_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_390/merge_stmt_403_PhiAck/dummy
      -- 
    if_choice_transition_1159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_397_branch_ack_1, ack => sendB_CP_1116_elements(1)); -- 
    cr_1181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(1), ack => type_cast_424_inst_req_1); -- 
    rr_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(1), ack => type_cast_424_inst_req_0); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_390/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_390/if_stmt_397_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_390/if_stmt_397_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_390/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_390/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_1163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_397_branch_ack_0, ack => sendB_CP_1116_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_sample_completed_
      -- 
    ra_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_424_inst_ack_0, ack => sendB_CP_1116_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/type_cast_424_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438/$exit
      -- CP-element group 4: 	 branch_block_stmt_390/assign_stmt_409_to_assign_stmt_438__exit__
      -- CP-element group 4: 	 branch_block_stmt_390/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/phi_stmt_441/$entry
      -- CP-element group 4: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$entry
      -- 
    ca_1182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_424_inst_ack_1, ack => sendB_CP_1116_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Sample/ack
      -- 
    ack_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_453_index_offset_ack_0, ack => sendB_CP_1116_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_request/req
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Update/$exit
      -- 
    ack_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_453_index_offset_ack_1, ack => sendB_CP_1116_elements(6)); -- 
    req_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(6), ack => addr_of_454_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_request/ack
      -- CP-element group 7: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_sample_completed_
      -- 
    ack_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_454_final_reg_ack_0, ack => sendB_CP_1116_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/word_access_start/word_0/rr
      -- 
    ack_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_454_final_reg_ack_1, ack => sendB_CP_1116_elements(8)); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(8), ack => ptr_deref_458_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Sample/word_access_start/word_0/ra
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_458_load_0_ack_0, ack => sendB_CP_1116_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	30 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/ptr_deref_458_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/ptr_deref_458_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/ptr_deref_458_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/ptr_deref_458_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Sample/rr
      -- 
    ca_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_458_load_0_ack_1, ack => sendB_CP_1116_elements(10)); -- 
    rr_1289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_504_inst_req_0); -- 
    rr_1317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_511_inst_req_0); -- 
    rr_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_518_inst_req_0); -- 
    rr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_525_inst_req_0); -- 
    rr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_532_inst_req_0); -- 
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_539_inst_req_0); -- 
    rr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_546_inst_req_0); -- 
    rr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(10), ack => type_cast_553_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Sample/ra
      -- 
    ra_1290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_0, ack => sendB_CP_1116_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Sample/req
      -- CP-element group 12: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Update/ca
      -- 
    ca_1295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_1, ack => sendB_CP_1116_elements(12)); -- 
    req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(12), ack => WPIPE_maxpool_output_pipe_506_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Update/req
      -- CP-element group 13: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Sample/ack
      -- CP-element group 13: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_update_start_
      -- 
    ack_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_506_inst_ack_0, ack => sendB_CP_1116_elements(13)); -- 
    req_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(13), ack => WPIPE_maxpool_output_pipe_506_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Update/ack
      -- CP-element group 14: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_506_Update/$exit
      -- 
    ack_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_506_inst_ack_1, ack => sendB_CP_1116_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_sample_completed_
      -- 
    ra_1318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_511_inst_ack_0, ack => sendB_CP_1116_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Update/ca
      -- 
    ca_1323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_511_inst_ack_1, ack => sendB_CP_1116_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Sample/req
      -- 
    req_1331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(17), ack => WPIPE_maxpool_output_pipe_513_inst_req_0); -- 
    sendB_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(14) & sendB_CP_1116_elements(16);
      gj_sendB_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_update_start_
      -- CP-element group 18: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Update/req
      -- 
    ack_1332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_513_inst_ack_0, ack => sendB_CP_1116_elements(18)); -- 
    req_1336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(18), ack => WPIPE_maxpool_output_pipe_513_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_513_Update/ack
      -- 
    ack_1337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_513_inst_ack_1, ack => sendB_CP_1116_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Sample/ra
      -- 
    ra_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_0, ack => sendB_CP_1116_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	58 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Update/ca
      -- 
    ca_1351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_1, ack => sendB_CP_1116_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Sample/req
      -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(22), ack => WPIPE_maxpool_output_pipe_520_inst_req_0); -- 
    sendB_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(19) & sendB_CP_1116_elements(21);
      gj_sendB_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_update_start_
      -- CP-element group 23: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Sample/ack
      -- CP-element group 23: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Update/req
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_520_inst_ack_0, ack => sendB_CP_1116_elements(23)); -- 
    req_1364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(23), ack => WPIPE_maxpool_output_pipe_520_inst_req_1); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_520_Update/ack
      -- 
    ack_1365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_520_inst_ack_1, ack => sendB_CP_1116_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Sample/ra
      -- 
    ra_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_0, ack => sendB_CP_1116_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Update/ca
      -- 
    ca_1379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_1, ack => sendB_CP_1116_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Sample/req
      -- 
    req_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(27), ack => WPIPE_maxpool_output_pipe_527_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(24) & sendB_CP_1116_elements(26);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_update_start_
      -- CP-element group 28: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Update/req
      -- 
    ack_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_527_inst_ack_0, ack => sendB_CP_1116_elements(28)); -- 
    req_1392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(28), ack => WPIPE_maxpool_output_pipe_527_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_527_Update/ack
      -- 
    ack_1393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_527_inst_ack_1, ack => sendB_CP_1116_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	10 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Sample/ra
      -- 
    ra_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_532_inst_ack_0, ack => sendB_CP_1116_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	58 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Update/ca
      -- 
    ca_1407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_532_inst_ack_1, ack => sendB_CP_1116_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Sample/req
      -- 
    req_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(32), ack => WPIPE_maxpool_output_pipe_534_inst_req_0); -- 
    sendB_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(29) & sendB_CP_1116_elements(31);
      gj_sendB_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_update_start_
      -- CP-element group 33: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Update/req
      -- 
    ack_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_534_inst_ack_0, ack => sendB_CP_1116_elements(33)); -- 
    req_1420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(33), ack => WPIPE_maxpool_output_pipe_534_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_534_Update/ack
      -- 
    ack_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_534_inst_ack_1, ack => sendB_CP_1116_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Sample/ra
      -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_0, ack => sendB_CP_1116_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	58 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Update/ca
      -- 
    ca_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_1, ack => sendB_CP_1116_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Sample/req
      -- 
    req_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(37), ack => WPIPE_maxpool_output_pipe_541_inst_req_0); -- 
    sendB_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(34) & sendB_CP_1116_elements(36);
      gj_sendB_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_update_start_
      -- CP-element group 38: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Update/req
      -- 
    ack_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_541_inst_ack_0, ack => sendB_CP_1116_elements(38)); -- 
    req_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(38), ack => WPIPE_maxpool_output_pipe_541_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_541_Update/ack
      -- 
    ack_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_541_inst_ack_1, ack => sendB_CP_1116_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Sample/ra
      -- 
    ra_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_546_inst_ack_0, ack => sendB_CP_1116_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Update/ca
      -- 
    ca_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_546_inst_ack_1, ack => sendB_CP_1116_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Sample/req
      -- 
    req_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(42), ack => WPIPE_maxpool_output_pipe_548_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(39) & sendB_CP_1116_elements(41);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_update_start_
      -- CP-element group 43: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Update/req
      -- 
    ack_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_548_inst_ack_0, ack => sendB_CP_1116_elements(43)); -- 
    req_1476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(43), ack => WPIPE_maxpool_output_pipe_548_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_548_Update/ack
      -- 
    ack_1477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_548_inst_ack_1, ack => sendB_CP_1116_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Sample/ra
      -- 
    ra_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_553_inst_ack_0, ack => sendB_CP_1116_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	58 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Update/ca
      -- 
    ca_1491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_553_inst_ack_1, ack => sendB_CP_1116_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Sample/req
      -- 
    req_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(47), ack => WPIPE_maxpool_output_pipe_555_inst_req_0); -- 
    sendB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(44) & sendB_CP_1116_elements(46);
      gj_sendB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_update_start_
      -- CP-element group 48: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Update/req
      -- 
    ack_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_555_inst_ack_0, ack => sendB_CP_1116_elements(48)); -- 
    req_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(48), ack => WPIPE_maxpool_output_pipe_555_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/WPIPE_maxpool_output_pipe_555_Update/ack
      -- 
    ack_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_555_inst_ack_1, ack => sendB_CP_1116_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/$exit
      -- CP-element group 50: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568__exit__
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569__entry__
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_390/R_exitcond1_570_place
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_390/if_stmt_569_else_link/$entry
      -- 
    branch_req_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(50), ack => if_stmt_569_branch_req_0); -- 
    sendB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(5) & sendB_CP_1116_elements(49);
      gj_sendB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_390/merge_stmt_575__exit__
      -- CP-element group 51: 	 branch_block_stmt_390/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_390/if_stmt_569_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_390/if_stmt_569_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_390/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_390/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_390/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_390/merge_stmt_575_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_390/merge_stmt_575_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_390/merge_stmt_575_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_390/merge_stmt_575_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_390/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_390/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_569_branch_ack_1, ack => sendB_CP_1116_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_390/if_stmt_569_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_390/if_stmt_569_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_569_branch_ack_0, ack => sendB_CP_1116_elements(52)); -- 
    rr_1566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(52), ack => type_cast_447_inst_req_0); -- 
    cr_1571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(52), ack => type_cast_447_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/phi_stmt_441/$exit
      -- CP-element group 53: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_445_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_390/bbx_xnph_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_req
      -- 
    phi_stmt_441_req_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_441_req_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(53), ack => phi_stmt_441_req_0); -- 
    -- Element group sendB_CP_1116_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendB_CP_1116_elements(4), ack => sendB_CP_1116_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/ra
      -- 
    ra_1567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_447_inst_ack_0, ack => sendB_CP_1116_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/ca
      -- 
    ca_1572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_447_inst_ack_1, ack => sendB_CP_1116_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/$exit
      -- CP-element group 56: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/$exit
      -- CP-element group 56: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_390/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_req
      -- 
    phi_stmt_441_req_1573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_441_req_1573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(56), ack => phi_stmt_441_req_1); -- 
    sendB_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1116_elements(54) & sendB_CP_1116_elements(55);
      gj_sendB_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1116_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_390/merge_stmt_440_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_390/merge_stmt_440_PhiAck/$entry
      -- 
    sendB_CP_1116_elements(57) <= OrReduce(sendB_CP_1116_elements(53) & sendB_CP_1116_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	21 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	31 
    -- CP-element group 58: 	36 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	46 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_complete/req
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/addr_of_454_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_504_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/ptr_deref_458_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_511_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/array_obj_ref_453_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/merge_stmt_440__exit__
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568__entry__
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_518_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_525_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_532_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_539_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_546_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_update_start_
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_390/assign_stmt_455_to_assign_stmt_568/type_cast_553_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_390/merge_stmt_440_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_390/merge_stmt_440_PhiAck/phi_stmt_441_ack
      -- 
    phi_stmt_441_ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_441_ack_0, ack => sendB_CP_1116_elements(58)); -- 
    cr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => ptr_deref_458_load_0_req_1); -- 
    req_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => addr_of_454_final_reg_req_1); -- 
    cr_1322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_511_inst_req_1); -- 
    req_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => array_obj_ref_453_index_offset_req_1); -- 
    req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => array_obj_ref_453_index_offset_req_0); -- 
    cr_1294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_504_inst_req_1); -- 
    cr_1350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_518_inst_req_1); -- 
    cr_1378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_525_inst_req_1); -- 
    cr_1406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_532_inst_req_1); -- 
    cr_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_539_inst_req_1); -- 
    cr_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_546_inst_req_1); -- 
    cr_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1116_elements(58), ack => type_cast_553_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_577__exit__
      -- CP-element group 59: 	 branch_block_stmt_390/return__
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_579__exit__
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_390/$exit
      -- CP-element group 59: 	 branch_block_stmt_390/branch_block_stmt_390__exit__
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_577_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_577_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_577_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_577_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_390/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_390/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_579_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_579_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_579_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_390/merge_stmt_579_PhiAck/dummy
      -- 
    sendB_CP_1116_elements(59) <= OrReduce(sendB_CP_1116_elements(2) & sendB_CP_1116_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_452_resized : std_logic_vector(13 downto 0);
    signal R_indvar_452_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_455 : std_logic_vector(31 downto 0);
    signal cmp76_396 : std_logic_vector(0 downto 0);
    signal conv52_505 : std_logic_vector(7 downto 0);
    signal conv55_512 : std_logic_vector(7 downto 0);
    signal conv58_519 : std_logic_vector(7 downto 0);
    signal conv61_526 : std_logic_vector(7 downto 0);
    signal conv64_533 : std_logic_vector(7 downto 0);
    signal conv67_540 : std_logic_vector(7 downto 0);
    signal conv70_547 : std_logic_vector(7 downto 0);
    signal conv73_554 : std_logic_vector(7 downto 0);
    signal exitcond1_568 : std_logic_vector(0 downto 0);
    signal iNsTr_1_425 : std_logic_vector(63 downto 0);
    signal indvar_441 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_563 : std_logic_vector(63 downto 0);
    signal ptr_deref_458_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_458_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_458_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_458_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_458_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_471 : std_logic_vector(63 downto 0);
    signal shr21_477 : std_logic_vector(63 downto 0);
    signal shr27_483 : std_logic_vector(63 downto 0);
    signal shr33_489 : std_logic_vector(63 downto 0);
    signal shr39_495 : std_logic_vector(63 downto 0);
    signal shr45_501 : std_logic_vector(63 downto 0);
    signal shr9_465 : std_logic_vector(63 downto 0);
    signal shr_409 : std_logic_vector(31 downto 0);
    signal shrx_xop_421 : std_logic_vector(31 downto 0);
    signal tmp4_459 : std_logic_vector(63 downto 0);
    signal tmp80_438 : std_logic_vector(63 downto 0);
    signal tmp_415 : std_logic_vector(0 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_407_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_413_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_429_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_445_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_447_wire : std_logic_vector(63 downto 0);
    signal type_cast_463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_469_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_475_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_481_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_487_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_561_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_431 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_453_constant_part_of_offset <= "00000000000000";
    array_obj_ref_453_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_453_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_453_resized_base_address <= "00000000000000";
    ptr_deref_458_word_offset_0 <= "00000000000000";
    type_cast_394_wire_constant <= "00000000000000000000000000000011";
    type_cast_407_wire_constant <= "00000000000000000000000000000010";
    type_cast_413_wire_constant <= "00000000000000000000000000000001";
    type_cast_419_wire_constant <= "11111111111111111111111111111111";
    type_cast_429_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_445_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_475_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_481_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_487_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_493_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_561_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_441: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_445_wire_constant & type_cast_447_wire;
      req <= phi_stmt_441_req_0 & phi_stmt_441_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_441",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_441_ack_0,
          idata => idata,
          odata => indvar_441,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_441
    -- flow-through select operator MUX_437_inst
    tmp80_438 <= xx_xop_431 when (tmp_415(0) /=  '0') else type_cast_436_wire_constant;
    addr_of_454_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_454_final_reg_req_0;
      addr_of_454_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_454_final_reg_req_1;
      addr_of_454_final_reg_ack_1<= rack(0);
      addr_of_454_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_454_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_453_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_424_inst_req_0;
      type_cast_424_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_424_inst_req_1;
      type_cast_424_inst_ack_1<= rack(0);
      type_cast_424_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_424_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xop_421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_1_425,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_447_inst_req_0;
      type_cast_447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_447_inst_req_1;
      type_cast_447_inst_ack_1<= rack(0);
      type_cast_447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_563,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_447_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_504_inst_req_0;
      type_cast_504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_504_inst_req_1;
      type_cast_504_inst_ack_1<= rack(0);
      type_cast_504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_511_inst_req_0;
      type_cast_511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_511_inst_req_1;
      type_cast_511_inst_ack_1<= rack(0);
      type_cast_511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_518_inst_req_0;
      type_cast_518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_518_inst_req_1;
      type_cast_518_inst_ack_1<= rack(0);
      type_cast_518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_525_inst_req_0;
      type_cast_525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_525_inst_req_1;
      type_cast_525_inst_ack_1<= rack(0);
      type_cast_525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_532_inst_req_0;
      type_cast_532_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_532_inst_req_1;
      type_cast_532_inst_ack_1<= rack(0);
      type_cast_532_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_532_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_477,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_533,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_539_inst_req_0;
      type_cast_539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_539_inst_req_1;
      type_cast_539_inst_ack_1<= rack(0);
      type_cast_539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_471,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_546_inst_req_0;
      type_cast_546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_546_inst_req_1;
      type_cast_546_inst_ack_1<= rack(0);
      type_cast_546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_553_inst_req_0;
      type_cast_553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_553_inst_req_1;
      type_cast_553_inst_ack_1<= rack(0);
      type_cast_553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_453_index_1_rename
    process(R_indvar_452_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_452_resized;
      ov(13 downto 0) := iv;
      R_indvar_452_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_453_index_1_resize
    process(indvar_441) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_441;
      ov := iv(13 downto 0);
      R_indvar_452_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_453_root_address_inst
    process(array_obj_ref_453_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_453_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_453_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_458_addr_0
    process(ptr_deref_458_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_458_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_458_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_458_base_resize
    process(arrayidx_455) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_455;
      ov := iv(13 downto 0);
      ptr_deref_458_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_458_gather_scatter
    process(ptr_deref_458_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_458_data_0;
      ov(63 downto 0) := iv;
      tmp4_459 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_458_root_address_inst
    process(ptr_deref_458_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_458_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_458_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_397_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp76_396;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_397_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_397_branch_req_0,
          ack0 => if_stmt_397_branch_ack_0,
          ack1 => if_stmt_397_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_569_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_568;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_569_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_569_branch_req_0,
          ack0 => if_stmt_569_branch_ack_0,
          ack1 => if_stmt_569_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_420_inst
    process(shr_409) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_409, type_cast_419_wire_constant, tmp_var);
      shrx_xop_421 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_430_inst
    process(iNsTr_1_425) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_425, type_cast_429_wire_constant, tmp_var);
      xx_xop_431 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_562_inst
    process(indvar_441) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_441, type_cast_561_wire_constant, tmp_var);
      indvarx_xnext_563 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_567_inst
    process(indvarx_xnext_563, tmp80_438) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_563, tmp80_438, tmp_var);
      exitcond1_568 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_408_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_407_wire_constant, tmp_var);
      shr_409 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_464_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_463_wire_constant, tmp_var);
      shr9_465 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_470_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_469_wire_constant, tmp_var);
      shr15_471 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_476_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_475_wire_constant, tmp_var);
      shr21_477 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_482_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_481_wire_constant, tmp_var);
      shr27_483 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_488_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_487_wire_constant, tmp_var);
      shr33_489 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_494_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_493_wire_constant, tmp_var);
      shr39_495 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_500_inst
    process(tmp4_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_459, type_cast_499_wire_constant, tmp_var);
      shr45_501 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_395_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_394_wire_constant, tmp_var);
      cmp76_396 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_414_inst
    process(shr_409) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_409, type_cast_413_wire_constant, tmp_var);
      tmp_415 <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_453_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_452_scaled;
      array_obj_ref_453_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_453_index_offset_req_0;
      array_obj_ref_453_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_453_index_offset_req_1;
      array_obj_ref_453_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_458_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_458_load_0_req_0;
      ptr_deref_458_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_458_load_0_req_1;
      ptr_deref_458_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_458_word_address_0;
      ptr_deref_458_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_506_inst WPIPE_maxpool_output_pipe_513_inst WPIPE_maxpool_output_pipe_520_inst WPIPE_maxpool_output_pipe_527_inst WPIPE_maxpool_output_pipe_534_inst WPIPE_maxpool_output_pipe_541_inst WPIPE_maxpool_output_pipe_548_inst WPIPE_maxpool_output_pipe_555_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_506_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_513_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_520_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_527_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_534_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_541_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_548_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_555_inst_req_0;
      WPIPE_maxpool_output_pipe_506_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_513_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_520_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_527_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_534_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_541_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_548_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_555_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_506_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_513_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_520_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_527_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_534_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_541_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_548_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_555_inst_req_1;
      WPIPE_maxpool_output_pipe_506_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_513_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_520_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_527_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_534_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_541_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_548_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_555_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv52_505 & conv55_512 & conv58_519 & conv61_526 & conv64_533 & conv67_540 & conv70_547 & conv73_554;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_307_start: Boolean;
  signal timer_CP_307_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_79_load_0_req_0 : boolean;
  signal LOAD_count_79_load_0_ack_0 : boolean;
  signal LOAD_count_79_load_0_req_1 : boolean;
  signal LOAD_count_79_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_307_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_307_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_307_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_307_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_307: Block -- control-path 
    signal timer_CP_307_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_307_elements(0) <= timer_CP_307_start;
    timer_CP_307_symbol <= timer_CP_307_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_80/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_sample_start_
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_update_start_
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Update/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_80/LOAD_count_79_Update/word_access_complete/word_0/cr
      -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_307_elements(0), ack => LOAD_count_79_load_0_req_1); -- 
    rr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_307_elements(0), ack => LOAD_count_79_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_80/LOAD_count_79_sample_completed_
      -- CP-element group 1: 	 assign_stmt_80/LOAD_count_79_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_80/LOAD_count_79_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_80/LOAD_count_79_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_80/LOAD_count_79_Sample/word_access_start/word_0/ra
      -- 
    ra_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_79_load_0_ack_0, ack => timer_CP_307_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_80/$exit
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_update_completed_
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/$exit
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/LOAD_count_79_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/LOAD_count_79_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/LOAD_count_79_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_80/LOAD_count_79_Update/LOAD_count_79_Merge/merge_ack
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_79_load_0_ack_1, ack => timer_CP_307_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_79_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_79_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_79_word_address_0 <= "0";
    -- equivalence LOAD_count_79_gather_scatter
    process(LOAD_count_79_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_79_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_79_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_79_load_0_req_0;
      LOAD_count_79_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_79_load_0_req_1;
      LOAD_count_79_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_79_word_address_0;
      LOAD_count_79_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_2656_start: Boolean;
  signal timerDaemon_CP_2656_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1107_branch_req_0 : boolean;
  signal phi_stmt_1109_req_1 : boolean;
  signal phi_stmt_1109_req_0 : boolean;
  signal phi_stmt_1109_ack_0 : boolean;
  signal ADD_u64_u64_1115_inst_req_0 : boolean;
  signal ADD_u64_u64_1115_inst_ack_0 : boolean;
  signal ADD_u64_u64_1115_inst_req_1 : boolean;
  signal ADD_u64_u64_1115_inst_ack_1 : boolean;
  signal STORE_count_1117_store_0_req_0 : boolean;
  signal STORE_count_1117_store_0_ack_0 : boolean;
  signal STORE_count_1117_store_0_req_1 : boolean;
  signal STORE_count_1117_store_0_ack_1 : boolean;
  signal do_while_stmt_1107_branch_ack_0 : boolean;
  signal do_while_stmt_1107_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_2656_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2656_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_2656_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2656_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_2656: Block -- control-path 
    signal timerDaemon_CP_2656_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_2656_elements(0) <= timerDaemon_CP_2656_start;
    timerDaemon_CP_2656_symbol <= timerDaemon_CP_2656_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1106/$entry
      -- CP-element group 0: 	 branch_block_stmt_1106/branch_block_stmt_1106__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1106/do_while_stmt_1107__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1106/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1106/branch_block_stmt_1106__exit__
      -- CP-element group 1: 	 branch_block_stmt_1106/do_while_stmt_1107__exit__
      -- 
    timerDaemon_CP_2656_elements(1) <= timerDaemon_CP_2656_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1106/do_while_stmt_1107/$entry
      -- CP-element group 2: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107__entry__
      -- 
    timerDaemon_CP_2656_elements(2) <= timerDaemon_CP_2656_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107__exit__
      -- 
    -- Element group timerDaemon_CP_2656_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_back
      -- 
    -- Element group timerDaemon_CP_2656_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1106/do_while_stmt_1107/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_taken/$entry
      -- 
    timerDaemon_CP_2656_elements(5) <= timerDaemon_CP_2656_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_body_done
      -- 
    timerDaemon_CP_2656_elements(6) <= timerDaemon_CP_2656_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_2656_elements(7) <= timerDaemon_CP_2656_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_2656_elements(8) <= timerDaemon_CP_2656_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_2656_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/condition_evaluated
      -- 
    condition_evaluated_2680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(10), ack => do_while_stmt_1107_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(35) & timerDaemon_CP_2656_elements(15);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(12) & timerDaemon_CP_2656_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(9) & timerDaemon_CP_2656_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(9) & timerDaemon_CP_2656_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_2656_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/aggregated_phi_update_ack
      -- 
    -- Element group timerDaemon_CP_2656_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_loopback_trigger
      -- 
    timerDaemon_CP_2656_elements(16) <= timerDaemon_CP_2656_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_loopback_sample_req_ps
      -- 
    phi_stmt_1109_loopback_sample_req_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1109_loopback_sample_req_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(17), ack => phi_stmt_1109_req_1); -- 
    -- Element group timerDaemon_CP_2656_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_entry_trigger
      -- 
    timerDaemon_CP_2656_elements(18) <= timerDaemon_CP_2656_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_entry_sample_req_ps
      -- CP-element group 19: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_entry_sample_req
      -- 
    phi_stmt_1109_entry_sample_req_2698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1109_entry_sample_req_2698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(19), ack => phi_stmt_1109_req_0); -- 
    -- Element group timerDaemon_CP_2656_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/phi_stmt_1109_phi_mux_ack_ps
      -- 
    phi_stmt_1109_phi_mux_ack_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1109_ack_0, ack => timerDaemon_CP_2656_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_sample_completed_
      -- 
    -- Element group timerDaemon_CP_2656_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_update_start_
      -- 
    -- Element group timerDaemon_CP_2656_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_update_completed__ps
      -- 
    timerDaemon_CP_2656_elements(23) <= timerDaemon_CP_2656_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/type_cast_1112_update_completed_
      -- 
    -- Element group timerDaemon_CP_2656_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_2656_elements(22), ack => timerDaemon_CP_2656_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_2656_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_update_start__ps
      -- 
    -- Element group timerDaemon_CP_2656_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Sample/rr
      -- 
    rr_2722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(27), ack => ADD_u64_u64_1115_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(25) & timerDaemon_CP_2656_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Update/cr
      -- 
    cr_2727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(28), ack => ADD_u64_u64_1115_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(26) & timerDaemon_CP_2656_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Sample/ra
      -- 
    ra_2723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1115_inst_ack_0, ack => timerDaemon_CP_2656_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/ADD_u64_u64_1115_Update/ca
      -- 
    ca_2728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1115_inst_ack_1, ack => timerDaemon_CP_2656_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/STORE_count_1117_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/STORE_count_1117_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/STORE_count_1117_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/STORE_count_1117_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/word_access_start/word_0/rr
      -- 
    rr_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(31), ack => STORE_count_1117_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(9) & timerDaemon_CP_2656_elements(15) & timerDaemon_CP_2656_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/word_access_complete/word_0/cr
      -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2656_elements(32), ack => STORE_count_1117_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_2656_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Sample/word_access_start/word_0/ra
      -- 
    ra_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1117_store_0_ack_0, ack => timerDaemon_CP_2656_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/STORE_count_1117_Update/word_access_complete/word_0/ca
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1117_store_0_ack_1, ack => timerDaemon_CP_2656_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_2656_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_2656_elements(9), ack => timerDaemon_CP_2656_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1106/do_while_stmt_1107/do_while_stmt_1107_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2656_elements(34) & timerDaemon_CP_2656_elements(14);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2656_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_exit/ack
      -- 
    ack_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1107_branch_ack_0, ack => timerDaemon_CP_2656_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_1106/do_while_stmt_1107/loop_taken/ack
      -- 
    ack_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1107_branch_ack_1, ack => timerDaemon_CP_2656_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1106/do_while_stmt_1107/$exit
      -- 
    timerDaemon_CP_2656_elements(39) <= timerDaemon_CP_2656_elements(3);
    timerDaemon_do_while_stmt_1107_terminator_2772: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1107_terminator_2772", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_2656_elements(6),loop_continue => timerDaemon_CP_2656_elements(38),loop_terminate => timerDaemon_CP_2656_elements(37),loop_back => timerDaemon_CP_2656_elements(4),loop_exit => timerDaemon_CP_2656_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1109_phi_seq_2729_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_2656_elements(18);
      timerDaemon_CP_2656_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_2656_elements(21);
      timerDaemon_CP_2656_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_2656_elements(23);
      timerDaemon_CP_2656_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_2656_elements(16);
      timerDaemon_CP_2656_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_2656_elements(29);
      timerDaemon_CP_2656_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_2656_elements(30);
      timerDaemon_CP_2656_elements(17) <= phi_mux_reqs(1);
      phi_stmt_1109_phi_seq_2729 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_1109_phi_seq_2729") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_2656_elements(11), 
          phi_sample_ack => timerDaemon_CP_2656_elements(14), 
          phi_update_req => timerDaemon_CP_2656_elements(13), 
          phi_update_ack => timerDaemon_CP_2656_elements(15), 
          phi_mux_ack => timerDaemon_CP_2656_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2681_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_2656_elements(7);
        preds(1)  <= timerDaemon_CP_2656_elements(8);
        entry_tmerge_2681 : transition_merge -- 
          generic map(name => " entry_tmerge_2681")
          port map (preds => preds, symbol_out => timerDaemon_CP_2656_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_1115_wire : std_logic_vector(63 downto 0);
    signal STORE_count_1117_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_1117_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_1114_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1121_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_1109 : std_logic_vector(63 downto 0);
    signal type_cast_1112_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_1117_word_address_0 <= "0";
    konst_1114_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1121_wire_constant <= "1";
    type_cast_1112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1109: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1112_wire_constant & ADD_u64_u64_1115_wire;
      req <= phi_stmt_1109_req_0 & phi_stmt_1109_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1109",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1109_ack_0,
          idata => idata,
          odata => ncount_1109,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1109
    -- equivalence STORE_count_1117_gather_scatter
    process(ncount_1109) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_1109;
      ov(63 downto 0) := iv;
      STORE_count_1117_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_1107_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1121_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1107_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1107_branch_req_0,
          ack0 => do_while_stmt_1107_branch_ack_0,
          ack1 => do_while_stmt_1107_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_1115_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_1109;
      ADD_u64_u64_1115_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1115_inst_req_0;
      ADD_u64_u64_1115_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1115_inst_req_1;
      ADD_u64_u64_1115_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_1117_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_1117_store_0_req_0;
      STORE_count_1117_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_1117_store_0_req_1;
      STORE_count_1117_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_1117_word_address_0;
      data_in <= STORE_count_1117_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module fill_T
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_T
  signal fill_T_addr :  std_logic_vector(63 downto 0);
  signal fill_T_in_args    : std_logic_vector(63 downto 0);
  signal fill_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_T_tag_out   : std_logic_vector(1 downto 0);
  signal fill_T_start_req : std_logic;
  signal fill_T_start_ack : std_logic;
  signal fill_T_fin_req   : std_logic;
  signal fill_T_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_T
  signal fill_T_call_reqs: std_logic_vector(0 downto 0);
  signal fill_T_call_acks: std_logic_vector(0 downto 0);
  signal fill_T_return_reqs: std_logic_vector(0 downto 0);
  signal fill_T_return_acks: std_logic_vector(0 downto 0);
  signal fill_T_call_data: std_logic_vector(63 downto 0);
  signal fill_T_call_tag: std_logic_vector(0 downto 0);
  signal fill_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module maxPool3D
  component maxPool3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      fill_T_call_reqs : out  std_logic_vector(0 downto 0);
      fill_T_call_acks : in   std_logic_vector(0 downto 0);
      fill_T_call_data : out  std_logic_vector(63 downto 0);
      fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_T_return_reqs : out  std_logic_vector(0 downto 0);
      fill_T_return_acks : in   std_logic_vector(0 downto 0);
      fill_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_call_acks : in   std_logic_vector(0 downto 0);
      maxPool4_call_data : out  std_logic_vector(159 downto 0);
      maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
      maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_return_acks : in   std_logic_vector(0 downto 0);
      maxPool4_return_data : in   std_logic_vector(7 downto 0);
      maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(31 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool3D
  signal maxPool3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool3D_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool3D_start_req : std_logic;
  signal maxPool3D_start_ack : std_logic;
  signal maxPool3D_fin_req   : std_logic;
  signal maxPool3D_fin_ack : std_logic;
  -- declarations related to module maxPool4
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool4
  signal maxPool4_addr :  std_logic_vector(31 downto 0);
  signal maxPool4_addr1 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr2 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr3 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr4 :  std_logic_vector(31 downto 0);
  signal maxPool4_output :  std_logic_vector(7 downto 0);
  signal maxPool4_in_args    : std_logic_vector(159 downto 0);
  signal maxPool4_out_args   : std_logic_vector(7 downto 0);
  signal maxPool4_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool4_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool4_start_req : std_logic;
  signal maxPool4_start_ack : std_logic;
  signal maxPool4_fin_req   : std_logic;
  signal maxPool4_fin_ack : std_logic;
  -- caller side aggregated signals for module maxPool4
  signal maxPool4_call_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_call_acks: std_logic_vector(0 downto 0);
  signal maxPool4_return_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_return_acks: std_logic_vector(0 downto 0);
  signal maxPool4_call_data: std_logic_vector(159 downto 0);
  signal maxPool4_call_tag: std_logic_vector(0 downto 0);
  signal maxPool4_return_data: std_logic_vector(7 downto 0);
  signal maxPool4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(31 downto 0);
  signal sendB_in_args    : std_logic_vector(31 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(31 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module fill_T
  fill_T_addr <= fill_T_in_args(63 downto 0);
  -- call arbiter for module fill_T
  fill_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_T_call_reqs,
      call_acks => fill_T_call_acks,
      return_reqs => fill_T_return_reqs,
      return_acks => fill_T_return_acks,
      call_data  => fill_T_call_data,
      call_tag  => fill_T_call_tag,
      return_tag  => fill_T_return_tag,
      call_mtag => fill_T_tag_in,
      return_mtag => fill_T_tag_out,
      call_mreq => fill_T_start_req,
      call_mack => fill_T_start_ack,
      return_mreq => fill_T_fin_req,
      return_mack => fill_T_fin_ack,
      call_mdata => fill_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  fill_T_instance:fill_T-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => fill_T_addr,
      start_req => fill_T_start_req,
      start_ack => fill_T_start_ack,
      fin_req => fill_T_fin_req,
      fin_ack => fill_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(1 downto 1),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(1 downto 1),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(15 downto 8),
      tag_in => fill_T_tag_in,
      tag_out => fill_T_tag_out-- 
    ); -- 
  -- module maxPool3D
  maxPool3D_instance:maxPool3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => maxPool3D_start_req,
      start_ack => maxPool3D_start_ack,
      fin_req => maxPool3D_fin_req,
      fin_ack => maxPool3D_fin_ack,
      clk => clk,
      reset => reset,
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      fill_T_call_reqs => fill_T_call_reqs(0 downto 0),
      fill_T_call_acks => fill_T_call_acks(0 downto 0),
      fill_T_call_data => fill_T_call_data(63 downto 0),
      fill_T_call_tag => fill_T_call_tag(0 downto 0),
      fill_T_return_reqs => fill_T_return_reqs(0 downto 0),
      fill_T_return_acks => fill_T_return_acks(0 downto 0),
      fill_T_return_tag => fill_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      maxPool4_call_reqs => maxPool4_call_reqs(0 downto 0),
      maxPool4_call_acks => maxPool4_call_acks(0 downto 0),
      maxPool4_call_data => maxPool4_call_data(159 downto 0),
      maxPool4_call_tag => maxPool4_call_tag(0 downto 0),
      maxPool4_return_reqs => maxPool4_return_reqs(0 downto 0),
      maxPool4_return_acks => maxPool4_return_acks(0 downto 0),
      maxPool4_return_data => maxPool4_return_data(7 downto 0),
      maxPool4_return_tag => maxPool4_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(31 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => maxPool3D_tag_in,
      tag_out => maxPool3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  maxPool3D_tag_in <= (others => '0');
  maxPool3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => maxPool3D_start_req, start_ack => maxPool3D_start_ack,  fin_req => maxPool3D_fin_req,  fin_ack => maxPool3D_fin_ack);
  -- module maxPool4
  maxPool4_addr <= maxPool4_in_args(159 downto 128);
  maxPool4_addr1 <= maxPool4_in_args(127 downto 96);
  maxPool4_addr2 <= maxPool4_in_args(95 downto 64);
  maxPool4_addr3 <= maxPool4_in_args(63 downto 32);
  maxPool4_addr4 <= maxPool4_in_args(31 downto 0);
  maxPool4_out_args <= maxPool4_output ;
  -- call arbiter for module maxPool4
  maxPool4_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 160,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => maxPool4_call_reqs,
      call_acks => maxPool4_call_acks,
      return_reqs => maxPool4_return_reqs,
      return_acks => maxPool4_return_acks,
      call_data  => maxPool4_call_data,
      call_tag  => maxPool4_call_tag,
      return_tag  => maxPool4_return_tag,
      call_mtag => maxPool4_tag_in,
      return_mtag => maxPool4_tag_out,
      return_data =>maxPool4_return_data,
      call_mreq => maxPool4_start_req,
      call_mack => maxPool4_start_ack,
      return_mreq => maxPool4_fin_req,
      return_mack => maxPool4_fin_ack,
      call_mdata => maxPool4_in_args,
      return_mdata => maxPool4_out_args,
      clk => clk, 
      reset => reset --
    ); --
  maxPool4_instance:maxPool4-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => maxPool4_addr,
      addr1 => maxPool4_addr1,
      addr2 => maxPool4_addr2,
      addr3 => maxPool4_addr3,
      addr4 => maxPool4_addr4,
      output => maxPool4_output,
      start_req => maxPool4_start_req,
      start_ack => maxPool4_start_ack,
      fin_req => maxPool4_fin_req,
      fin_ack => maxPool4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => maxPool4_tag_in,
      tag_out => maxPool4_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(31 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
