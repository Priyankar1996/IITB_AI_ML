-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_34_start: Boolean;
  signal convTranspose_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_1055_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1102_inst_req_1 : boolean;
  signal type_cast_691_inst_req_0 : boolean;
  signal type_cast_691_inst_ack_0 : boolean;
  signal type_cast_471_inst_ack_1 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal type_cast_691_inst_req_1 : boolean;
  signal type_cast_691_inst_ack_1 : boolean;
  signal addr_of_671_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 : boolean;
  signal type_cast_471_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1090_inst_req_0 : boolean;
  signal type_cast_1075_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_480_inst_ack_1 : boolean;
  signal ptr_deref_600_store_0_req_0 : boolean;
  signal type_cast_502_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_480_inst_req_1 : boolean;
  signal type_cast_471_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_480_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_480_inst_req_0 : boolean;
  signal addr_of_671_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal if_stmt_1112_branch_ack_0 : boolean;
  signal ptr_deref_600_store_0_ack_0 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal type_cast_471_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_467_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal call_stmt_1002_call_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_674_inst_ack_1 : boolean;
  signal array_obj_ref_670_index_offset_ack_0 : boolean;
  signal type_cast_502_inst_req_1 : boolean;
  signal type_cast_1065_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_1015_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal if_stmt_614_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 : boolean;
  signal array_obj_ref_1168_index_offset_req_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_674_inst_req_1 : boolean;
  signal array_obj_ref_670_index_offset_req_0 : boolean;
  signal type_cast_556_inst_ack_1 : boolean;
  signal type_cast_502_inst_ack_0 : boolean;
  signal call_stmt_1002_call_req_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal addr_of_671_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_req_1 : boolean;
  signal type_cast_556_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal call_stmt_1002_call_req_0 : boolean;
  signal type_cast_101_inst_req_0 : boolean;
  signal type_cast_101_inst_ack_0 : boolean;
  signal type_cast_101_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 : boolean;
  signal type_cast_101_inst_ack_1 : boolean;
  signal addr_of_671_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_467_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal type_cast_502_inst_req_0 : boolean;
  signal type_cast_556_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_467_inst_req_1 : boolean;
  signal type_cast_574_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 : boolean;
  signal type_cast_556_inst_req_0 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1096_inst_req_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal type_cast_574_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_325_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_325_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_325_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_325_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_0 : boolean;
  signal type_cast_1065_inst_req_1 : boolean;
  signal type_cast_329_inst_req_0 : boolean;
  signal type_cast_329_inst_ack_0 : boolean;
  signal type_cast_329_inst_req_1 : boolean;
  signal type_cast_329_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_467_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_674_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal type_cast_574_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_674_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1108_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1087_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 : boolean;
  signal type_cast_1015_inst_req_0 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1102_inst_ack_1 : boolean;
  signal type_cast_641_inst_ack_1 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal type_cast_188_inst_req_0 : boolean;
  signal type_cast_188_inst_ack_0 : boolean;
  signal type_cast_188_inst_req_1 : boolean;
  signal type_cast_188_inst_ack_1 : boolean;
  signal type_cast_1139_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 : boolean;
  signal addr_of_464_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 : boolean;
  signal type_cast_641_inst_req_1 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_1015_inst_ack_1 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal type_cast_1015_inst_ack_0 : boolean;
  signal type_cast_210_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal type_cast_210_inst_ack_0 : boolean;
  signal type_cast_1006_inst_ack_1 : boolean;
  signal type_cast_210_inst_req_1 : boolean;
  signal type_cast_210_inst_ack_1 : boolean;
  signal type_cast_1139_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1087_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_1 : boolean;
  signal type_cast_218_inst_req_0 : boolean;
  signal type_cast_218_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1090_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal type_cast_218_inst_req_1 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_218_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 : boolean;
  signal call_stmt_1002_call_ack_1 : boolean;
  signal type_cast_232_inst_req_0 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_232_inst_ack_0 : boolean;
  signal type_cast_232_inst_req_1 : boolean;
  signal type_cast_232_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_0 : boolean;
  signal type_cast_908_inst_req_0 : boolean;
  signal type_cast_236_inst_req_0 : boolean;
  signal type_cast_236_inst_ack_0 : boolean;
  signal type_cast_236_inst_req_1 : boolean;
  signal type_cast_236_inst_ack_1 : boolean;
  signal type_cast_678_inst_ack_1 : boolean;
  signal type_cast_240_inst_req_0 : boolean;
  signal type_cast_240_inst_ack_0 : boolean;
  signal type_cast_240_inst_req_1 : boolean;
  signal type_cast_240_inst_ack_1 : boolean;
  signal type_cast_678_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal type_cast_244_inst_req_0 : boolean;
  signal type_cast_244_inst_ack_0 : boolean;
  signal type_cast_244_inst_req_1 : boolean;
  signal type_cast_244_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal addr_of_464_final_reg_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1087_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1108_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_ack_1 : boolean;
  signal type_cast_641_inst_ack_0 : boolean;
  signal type_cast_1006_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal type_cast_266_inst_req_0 : boolean;
  signal type_cast_266_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_1 : boolean;
  signal type_cast_266_inst_ack_1 : boolean;
  signal ptr_deref_600_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_275_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_275_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_275_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_275_inst_ack_1 : boolean;
  signal type_cast_641_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_1 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal type_cast_279_inst_req_0 : boolean;
  signal type_cast_279_inst_ack_0 : boolean;
  signal type_cast_279_inst_req_1 : boolean;
  signal type_cast_279_inst_ack_1 : boolean;
  signal array_obj_ref_670_index_offset_ack_1 : boolean;
  signal ptr_deref_600_store_0_req_1 : boolean;
  signal type_cast_678_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_ack_0 : boolean;
  signal addr_of_464_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_ack_1 : boolean;
  signal type_cast_291_inst_req_0 : boolean;
  signal type_cast_291_inst_ack_0 : boolean;
  signal type_cast_291_inst_req_1 : boolean;
  signal type_cast_291_inst_ack_1 : boolean;
  signal type_cast_678_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1096_inst_ack_1 : boolean;
  signal addr_of_464_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_300_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_300_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_300_inst_req_1 : boolean;
  signal type_cast_1075_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_300_inst_ack_1 : boolean;
  signal type_cast_1075_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 : boolean;
  signal type_cast_304_inst_req_0 : boolean;
  signal type_cast_304_inst_ack_0 : boolean;
  signal type_cast_304_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_1 : boolean;
  signal type_cast_304_inst_ack_1 : boolean;
  signal array_obj_ref_670_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal type_cast_316_inst_req_0 : boolean;
  signal type_cast_316_inst_ack_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_1 : boolean;
  signal type_cast_316_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_ack_0 : boolean;
  signal array_obj_ref_463_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_ack_1 : boolean;
  signal type_cast_341_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1099_inst_req_0 : boolean;
  signal type_cast_341_inst_ack_0 : boolean;
  signal type_cast_1065_inst_ack_1 : boolean;
  signal type_cast_341_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_0 : boolean;
  signal type_cast_341_inst_ack_1 : boolean;
  signal array_obj_ref_463_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_350_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_350_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_350_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_350_inst_ack_1 : boolean;
  signal type_cast_1065_inst_req_0 : boolean;
  signal type_cast_484_inst_ack_1 : boolean;
  signal type_cast_484_inst_req_1 : boolean;
  signal type_cast_354_inst_req_0 : boolean;
  signal type_cast_354_inst_ack_0 : boolean;
  signal type_cast_354_inst_req_1 : boolean;
  signal type_cast_354_inst_ack_1 : boolean;
  signal array_obj_ref_463_index_offset_ack_0 : boolean;
  signal array_obj_ref_463_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_ack_1 : boolean;
  signal if_stmt_614_branch_ack_0 : boolean;
  signal type_cast_484_inst_ack_0 : boolean;
  signal type_cast_484_inst_req_0 : boolean;
  signal type_cast_366_inst_req_0 : boolean;
  signal type_cast_366_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1087_inst_ack_1 : boolean;
  signal type_cast_366_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1099_inst_ack_0 : boolean;
  signal type_cast_366_inst_ack_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal type_cast_1006_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_375_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_375_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_375_inst_req_1 : boolean;
  signal type_cast_1006_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_375_inst_ack_1 : boolean;
  signal if_stmt_614_branch_ack_1 : boolean;
  signal type_cast_379_inst_req_0 : boolean;
  signal type_cast_379_inst_ack_0 : boolean;
  signal type_cast_379_inst_req_1 : boolean;
  signal type_cast_379_inst_ack_1 : boolean;
  signal type_cast_1075_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1090_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1090_inst_ack_1 : boolean;
  signal if_stmt_392_branch_req_0 : boolean;
  signal WPIPE_Block0_start_993_inst_req_0 : boolean;
  signal if_stmt_392_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_0 : boolean;
  signal if_stmt_392_branch_ack_0 : boolean;
  signal if_stmt_407_branch_req_0 : boolean;
  signal if_stmt_407_branch_ack_1 : boolean;
  signal if_stmt_407_branch_ack_0 : boolean;
  signal type_cast_434_inst_req_0 : boolean;
  signal type_cast_434_inst_ack_0 : boolean;
  signal type_cast_434_inst_req_1 : boolean;
  signal type_cast_434_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1105_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 : boolean;
  signal type_cast_1139_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1096_inst_ack_0 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal array_obj_ref_1168_index_offset_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1102_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1105_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1096_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 : boolean;
  signal type_cast_1139_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1102_inst_req_0 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 : boolean;
  signal if_stmt_1112_branch_ack_1 : boolean;
  signal type_cast_745_inst_req_0 : boolean;
  signal type_cast_745_inst_ack_0 : boolean;
  signal type_cast_745_inst_req_1 : boolean;
  signal type_cast_745_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1105_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1105_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 : boolean;
  signal type_cast_1045_inst_ack_1 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal type_cast_763_inst_req_1 : boolean;
  signal type_cast_763_inst_ack_1 : boolean;
  signal array_obj_ref_1168_index_offset_ack_0 : boolean;
  signal RPIPE_Block0_done_998_inst_ack_1 : boolean;
  signal type_cast_1045_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_0 : boolean;
  signal type_cast_1162_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_998_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 : boolean;
  signal type_cast_1045_inst_ack_0 : boolean;
  signal type_cast_1045_inst_req_0 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_0 : boolean;
  signal type_cast_1162_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_998_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_998_inst_req_0 : boolean;
  signal if_stmt_1112_branch_req_0 : boolean;
  signal type_cast_908_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal type_cast_1035_inst_ack_1 : boolean;
  signal type_cast_1035_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1093_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1093_inst_req_1 : boolean;
  signal ptr_deref_807_store_0_req_0 : boolean;
  signal ptr_deref_807_store_0_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal ptr_deref_807_store_0_req_1 : boolean;
  signal ptr_deref_807_store_0_ack_1 : boolean;
  signal array_obj_ref_1168_index_offset_ack_1 : boolean;
  signal type_cast_1035_inst_ack_0 : boolean;
  signal type_cast_1035_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1108_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1108_inst_req_0 : boolean;
  signal if_stmt_821_branch_req_0 : boolean;
  signal if_stmt_821_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_1 : boolean;
  signal if_stmt_821_branch_ack_0 : boolean;
  signal type_cast_1085_inst_ack_1 : boolean;
  signal type_cast_832_inst_req_0 : boolean;
  signal type_cast_832_inst_ack_0 : boolean;
  signal type_cast_1085_inst_req_1 : boolean;
  signal type_cast_832_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1093_inst_ack_0 : boolean;
  signal type_cast_832_inst_ack_1 : boolean;
  signal type_cast_836_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1093_inst_req_0 : boolean;
  signal type_cast_836_inst_ack_0 : boolean;
  signal type_cast_836_inst_req_1 : boolean;
  signal type_cast_836_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1099_inst_ack_1 : boolean;
  signal type_cast_1025_inst_ack_1 : boolean;
  signal type_cast_1025_inst_req_1 : boolean;
  signal type_cast_840_inst_req_0 : boolean;
  signal type_cast_840_inst_ack_0 : boolean;
  signal type_cast_840_inst_req_1 : boolean;
  signal type_cast_840_inst_ack_1 : boolean;
  signal if_stmt_858_branch_req_0 : boolean;
  signal type_cast_1025_inst_ack_0 : boolean;
  signal if_stmt_858_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_983_inst_req_1 : boolean;
  signal if_stmt_858_branch_ack_0 : boolean;
  signal type_cast_1085_inst_ack_0 : boolean;
  signal type_cast_1085_inst_req_0 : boolean;
  signal type_cast_1025_inst_req_0 : boolean;
  signal type_cast_885_inst_req_0 : boolean;
  signal type_cast_885_inst_ack_0 : boolean;
  signal type_cast_885_inst_req_1 : boolean;
  signal type_cast_885_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1099_inst_req_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_1 : boolean;
  signal array_obj_ref_914_index_offset_req_0 : boolean;
  signal array_obj_ref_914_index_offset_ack_0 : boolean;
  signal array_obj_ref_914_index_offset_req_1 : boolean;
  signal array_obj_ref_914_index_offset_ack_1 : boolean;
  signal addr_of_915_final_reg_req_0 : boolean;
  signal addr_of_915_final_reg_ack_0 : boolean;
  signal addr_of_915_final_reg_req_1 : boolean;
  signal addr_of_915_final_reg_ack_1 : boolean;
  signal type_cast_1162_inst_req_1 : boolean;
  signal type_cast_1162_inst_ack_1 : boolean;
  signal ptr_deref_918_store_0_req_0 : boolean;
  signal ptr_deref_918_store_0_ack_0 : boolean;
  signal type_cast_908_inst_req_1 : boolean;
  signal ptr_deref_918_store_0_req_1 : boolean;
  signal ptr_deref_918_store_0_ack_1 : boolean;
  signal type_cast_908_inst_ack_1 : boolean;
  signal phi_stmt_1156_req_1 : boolean;
  signal if_stmt_933_branch_req_0 : boolean;
  signal phi_stmt_902_req_1 : boolean;
  signal if_stmt_933_branch_ack_1 : boolean;
  signal if_stmt_933_branch_ack_0 : boolean;
  signal call_stmt_944_call_req_0 : boolean;
  signal call_stmt_944_call_ack_0 : boolean;
  signal call_stmt_944_call_req_1 : boolean;
  signal call_stmt_944_call_ack_1 : boolean;
  signal type_cast_949_inst_req_0 : boolean;
  signal type_cast_949_inst_ack_0 : boolean;
  signal type_cast_949_inst_req_1 : boolean;
  signal type_cast_949_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_952_inst_req_0 : boolean;
  signal WPIPE_Block0_start_952_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_952_inst_req_1 : boolean;
  signal WPIPE_Block0_start_952_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_955_inst_req_0 : boolean;
  signal WPIPE_Block0_start_955_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_955_inst_req_1 : boolean;
  signal WPIPE_Block0_start_955_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_958_inst_req_0 : boolean;
  signal WPIPE_Block0_start_958_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_958_inst_req_1 : boolean;
  signal WPIPE_Block0_start_958_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_961_inst_req_0 : boolean;
  signal WPIPE_Block0_start_961_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_961_inst_req_1 : boolean;
  signal WPIPE_Block0_start_961_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_964_inst_req_0 : boolean;
  signal WPIPE_Block0_start_964_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_964_inst_req_1 : boolean;
  signal WPIPE_Block0_start_964_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_967_inst_req_0 : boolean;
  signal WPIPE_Block0_start_967_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_967_inst_req_1 : boolean;
  signal WPIPE_Block0_start_967_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_970_inst_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_1 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_973_inst_req_0 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_973_inst_req_1 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_976_inst_req_0 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_976_inst_req_1 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_979_inst_req_0 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_979_inst_req_1 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_983_inst_req_0 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_0 : boolean;
  signal addr_of_1169_final_reg_req_0 : boolean;
  signal addr_of_1169_final_reg_ack_0 : boolean;
  signal addr_of_1169_final_reg_req_1 : boolean;
  signal addr_of_1169_final_reg_ack_1 : boolean;
  signal ptr_deref_1173_load_0_req_0 : boolean;
  signal ptr_deref_1173_load_0_ack_0 : boolean;
  signal ptr_deref_1173_load_0_req_1 : boolean;
  signal ptr_deref_1173_load_0_ack_1 : boolean;
  signal type_cast_1177_inst_req_0 : boolean;
  signal type_cast_1177_inst_ack_0 : boolean;
  signal type_cast_1177_inst_req_1 : boolean;
  signal type_cast_1177_inst_ack_1 : boolean;
  signal type_cast_1187_inst_req_0 : boolean;
  signal type_cast_1187_inst_ack_0 : boolean;
  signal type_cast_1187_inst_req_1 : boolean;
  signal type_cast_1187_inst_ack_1 : boolean;
  signal type_cast_1197_inst_req_0 : boolean;
  signal type_cast_1197_inst_ack_0 : boolean;
  signal type_cast_1197_inst_req_1 : boolean;
  signal type_cast_1197_inst_ack_1 : boolean;
  signal type_cast_1207_inst_req_0 : boolean;
  signal type_cast_1207_inst_ack_0 : boolean;
  signal type_cast_1207_inst_req_1 : boolean;
  signal type_cast_1207_inst_ack_1 : boolean;
  signal type_cast_1217_inst_req_0 : boolean;
  signal type_cast_1217_inst_ack_0 : boolean;
  signal type_cast_1217_inst_req_1 : boolean;
  signal type_cast_1217_inst_ack_1 : boolean;
  signal type_cast_1227_inst_req_0 : boolean;
  signal type_cast_1227_inst_ack_0 : boolean;
  signal type_cast_1227_inst_req_1 : boolean;
  signal type_cast_1227_inst_ack_1 : boolean;
  signal type_cast_1237_inst_req_0 : boolean;
  signal type_cast_1237_inst_ack_0 : boolean;
  signal type_cast_1237_inst_req_1 : boolean;
  signal type_cast_1237_inst_ack_1 : boolean;
  signal type_cast_1247_inst_req_0 : boolean;
  signal type_cast_1247_inst_ack_0 : boolean;
  signal type_cast_1247_inst_req_1 : boolean;
  signal type_cast_1247_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_ack_0 : boolean;
  signal phi_stmt_1156_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_ack_1 : boolean;
  signal if_stmt_1284_branch_req_0 : boolean;
  signal phi_stmt_902_ack_0 : boolean;
  signal if_stmt_1284_branch_ack_1 : boolean;
  signal if_stmt_1284_branch_ack_0 : boolean;
  signal phi_stmt_451_req_0 : boolean;
  signal type_cast_457_inst_req_0 : boolean;
  signal type_cast_457_inst_ack_0 : boolean;
  signal type_cast_457_inst_req_1 : boolean;
  signal type_cast_457_inst_ack_1 : boolean;
  signal phi_stmt_451_req_1 : boolean;
  signal phi_stmt_451_ack_0 : boolean;
  signal phi_stmt_658_req_0 : boolean;
  signal type_cast_664_inst_req_0 : boolean;
  signal type_cast_664_inst_ack_0 : boolean;
  signal type_cast_664_inst_req_1 : boolean;
  signal type_cast_664_inst_ack_1 : boolean;
  signal phi_stmt_658_req_1 : boolean;
  signal phi_stmt_902_req_0 : boolean;
  signal phi_stmt_658_ack_0 : boolean;
  signal phi_stmt_1156_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_34: Block -- control-path 
    signal convTranspose_CP_34_elements: BooleanArray(387 downto 0);
    -- 
  begin -- 
    convTranspose_CP_34_elements(0) <= convTranspose_CP_34_start;
    convTranspose_CP_34_symbol <= convTranspose_CP_34_elements(387);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Update/cr
      -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_138_inst_req_1); -- 
    cr_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_51_inst_req_1); -- 
    cr_207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_76_inst_req_1); -- 
    cr_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_101_inst_req_1); -- 
    cr_319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_329_inst_req_1); -- 
    cr_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_163_inst_req_1); -- 
    cr_459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_188_inst_req_1); -- 
    cr_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_201_inst_req_1); -- 
    cr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_210_inst_req_1); -- 
    cr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_214_inst_req_1); -- 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_218_inst_req_1); -- 
    cr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_232_inst_req_1); -- 
    cr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_236_inst_req_1); -- 
    cr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_240_inst_req_1); -- 
    cr_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_244_inst_req_1); -- 
    cr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_266_inst_req_1); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_279_inst_req_1); -- 
    cr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_291_inst_req_1); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_304_inst_req_1); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_316_inst_req_1); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_341_inst_req_1); -- 
    cr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_354_inst_req_1); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_366_inst_req_1); -- 
    cr_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_379_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => convTranspose_CP_34_elements(1)); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Sample/rr
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => convTranspose_CP_34_elements(2)); -- 
    rr_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Sample/ra
      -- 
    ra_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => convTranspose_CP_34_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_38_Update/ca
      -- 
    ca_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => convTranspose_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_update_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Update/cr
      -- 
    ra_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_0, ack => convTranspose_CP_34_elements(5)); -- 
    cr_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(5), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_47_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_1, ack => convTranspose_CP_34_elements(6)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => type_cast_51_inst_req_0); -- 
    rr_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Sample/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => convTranspose_CP_34_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_51_Update/ca
      -- 
    ca_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => convTranspose_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => convTranspose_CP_34_elements(9)); -- 
    cr_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Sample/rr
      -- 
    ca_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => convTranspose_CP_34_elements(10)); -- 
    rr_202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => type_cast_63_inst_req_0); -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Sample/ra
      -- 
    ra_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => convTranspose_CP_34_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_63_Update/ca
      -- 
    ca_208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => convTranspose_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_update_start_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Update/cr
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_0, ack => convTranspose_CP_34_elements(13)); -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(13), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_72_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Sample/rr
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_1, ack => convTranspose_CP_34_elements(14)); -- 
    rr_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_0); -- 
    rr_230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => type_cast_76_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Sample/ra
      -- 
    ra_231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => convTranspose_CP_34_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_76_Update/ca
      -- 
    ca_236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => convTranspose_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_update_start_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Update/cr
      -- 
    ra_245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_0, ack => convTranspose_CP_34_elements(17)); -- 
    cr_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(17), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_84_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_1, ack => convTranspose_CP_34_elements(18)); -- 
    rr_258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => type_cast_88_inst_req_0); -- 
    rr_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Sample/ra
      -- 
    ra_259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => convTranspose_CP_34_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_88_Update/ca
      -- 
    ca_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => convTranspose_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_34_elements(21)); -- 
    cr_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(21), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Sample/rr
      -- 
    ca_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_34_elements(22)); -- 
    rr_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => type_cast_101_inst_req_0); -- 
    rr_300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Sample/ra
      -- 
    ra_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_0, ack => convTranspose_CP_34_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_101_Update/ca
      -- 
    ca_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_1, ack => convTranspose_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_update_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Update/cr
      -- 
    ra_301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_0, ack => convTranspose_CP_34_elements(25)); -- 
    cr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(25), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_109_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Sample/rr
      -- 
    ca_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_1, ack => convTranspose_CP_34_elements(26)); -- 
    rr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_0); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => type_cast_113_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Sample/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => convTranspose_CP_34_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_113_Update/ca
      -- 
    ca_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => convTranspose_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Update/cr
      -- 
    ra_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_0, ack => convTranspose_CP_34_elements(29)); -- 
    cr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(29), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_122_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Sample/rr
      -- 
    ca_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_1, ack => convTranspose_CP_34_elements(30)); -- 
    rr_342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => type_cast_126_inst_req_0); -- 
    rr_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Sample/ra
      -- 
    ra_343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => convTranspose_CP_34_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_126_Update/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => convTranspose_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_update_start_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Update/cr
      -- 
    ra_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_0, ack => convTranspose_CP_34_elements(33)); -- 
    cr_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(33), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_134_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Sample/rr
      -- 
    ca_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_1, ack => convTranspose_CP_34_elements(34)); -- 
    rr_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_0); -- 
    rr_370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => type_cast_138_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_sample_completed_
      -- 
    ra_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => convTranspose_CP_34_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_138_Update/ca
      -- 
    ca_376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => convTranspose_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_update_start_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Update/cr
      -- 
    ra_385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_0, ack => convTranspose_CP_34_elements(37)); -- 
    cr_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(37), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_147_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_1, ack => convTranspose_CP_34_elements(38)); -- 
    rr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    rr_398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => type_cast_151_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Sample/ra
      -- 
    ra_399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_34_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_151_Update/ca
      -- 
    ca_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_34_elements(41)); -- 
    cr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(41), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Sample/rr
      -- 
    ca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_34_elements(42)); -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_0); -- 
    rr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => type_cast_163_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Sample/ra
      -- 
    ra_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => convTranspose_CP_34_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_163_Update/ca
      -- 
    ca_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => convTranspose_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_update_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Update/cr
      -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_0, ack => convTranspose_CP_34_elements(45)); -- 
    cr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(45), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_172_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Sample/rr
      -- 
    ca_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_1, ack => convTranspose_CP_34_elements(46)); -- 
    rr_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => type_cast_176_inst_req_0); -- 
    rr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Sample/ra
      -- 
    ra_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => convTranspose_CP_34_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_176_Update/ca
      -- 
    ca_460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => convTranspose_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_update_start_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Update/cr
      -- 
    ra_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_0, ack => convTranspose_CP_34_elements(49)); -- 
    cr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(49), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_184_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Sample/rr
      -- 
    ca_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_1, ack => convTranspose_CP_34_elements(50)); -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => type_cast_188_inst_req_0); -- 
    rr_496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Sample/ra
      -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_0, ack => convTranspose_CP_34_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_188_Update/ca
      -- 
    ca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_1, ack => convTranspose_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_update_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Update/cr
      -- 
    ra_497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_0, ack => convTranspose_CP_34_elements(53)); -- 
    cr_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(53), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_197_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Sample/rr
      -- 
    ca_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_1, ack => convTranspose_CP_34_elements(54)); -- 
    rr_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => type_cast_201_inst_req_0); -- 
    rr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => RPIPE_ConvTranspose_input_pipe_262_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Sample/ra
      -- 
    ra_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => convTranspose_CP_34_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_201_Update/ca
      -- 
    ca_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => convTranspose_CP_34_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Sample/rr
      -- 
    rr_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(57), ack => type_cast_210_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(4) & convTranspose_CP_34_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Sample/ra
      -- 
    ra_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_0, ack => convTranspose_CP_34_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_210_Update/ca
      -- 
    ca_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_1, ack => convTranspose_CP_34_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	12 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Sample/rr
      -- 
    rr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(60), ack => type_cast_214_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(16) & convTranspose_CP_34_elements(12);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Sample/ra
      -- 
    ra_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => convTranspose_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_214_Update/ca
      -- 
    ca_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => convTranspose_CP_34_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	24 
    -- CP-element group 63: 	20 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Sample/rr
      -- 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(63), ack => type_cast_218_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(24) & convTranspose_CP_34_elements(20);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Sample/ra
      -- 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_0, ack => convTranspose_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_218_Update/ca
      -- 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_1, ack => convTranspose_CP_34_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	28 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Sample/rr
      -- 
    rr_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(66), ack => type_cast_232_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(32) & convTranspose_CP_34_elements(28);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Sample/ra
      -- 
    ra_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_232_inst_ack_0, ack => convTranspose_CP_34_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_232_Update/ca
      -- 
    ca_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_232_inst_ack_1, ack => convTranspose_CP_34_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Sample/rr
      -- 
    rr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(69), ack => type_cast_236_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(40) & convTranspose_CP_34_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Sample/ra
      -- 
    ra_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_236_inst_ack_0, ack => convTranspose_CP_34_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_236_Update/ca
      -- 
    ca_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_236_inst_ack_1, ack => convTranspose_CP_34_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Sample/rr
      -- 
    rr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(72), ack => type_cast_240_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(44) & convTranspose_CP_34_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Sample/ra
      -- 
    ra_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_240_inst_ack_0, ack => convTranspose_CP_34_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_240_Update/ca
      -- 
    ca_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_240_inst_ack_1, ack => convTranspose_CP_34_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Sample/rr
      -- 
    rr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(75), ack => type_cast_244_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(52) & convTranspose_CP_34_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Sample/ra
      -- 
    ra_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_244_inst_ack_0, ack => convTranspose_CP_34_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_244_Update/ca
      -- 
    ca_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_244_inst_ack_1, ack => convTranspose_CP_34_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_update_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Update/cr
      -- 
    ra_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_262_inst_ack_0, ack => convTranspose_CP_34_elements(78)); -- 
    cr_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(78), ack => RPIPE_ConvTranspose_input_pipe_262_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_262_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Sample/rr
      -- 
    ca_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_262_inst_ack_1, ack => convTranspose_CP_34_elements(79)); -- 
    rr_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => type_cast_266_inst_req_0); -- 
    rr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => RPIPE_ConvTranspose_input_pipe_275_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Sample/ra
      -- 
    ra_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_0, ack => convTranspose_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_266_Update/ca
      -- 
    ca_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_1, ack => convTranspose_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_update_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Update/cr
      -- 
    ra_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_275_inst_ack_0, ack => convTranspose_CP_34_elements(82)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(82), ack => RPIPE_ConvTranspose_input_pipe_275_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_275_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Sample/rr
      -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_275_inst_ack_1, ack => convTranspose_CP_34_elements(83)); -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => type_cast_279_inst_req_0); -- 
    rr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => RPIPE_ConvTranspose_input_pipe_287_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Sample/ra
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_279_inst_ack_0, ack => convTranspose_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_279_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_279_inst_ack_1, ack => convTranspose_CP_34_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_update_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Update/cr
      -- 
    ra_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_287_inst_ack_0, ack => convTranspose_CP_34_elements(86)); -- 
    cr_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(86), ack => RPIPE_ConvTranspose_input_pipe_287_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_287_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Sample/rr
      -- 
    ca_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_287_inst_ack_1, ack => convTranspose_CP_34_elements(87)); -- 
    rr_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => RPIPE_ConvTranspose_input_pipe_300_inst_req_0); -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => type_cast_291_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Sample/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_0, ack => convTranspose_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_291_Update/ca
      -- 
    ca_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_1, ack => convTranspose_CP_34_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Update/cr
      -- 
    ra_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_300_inst_ack_0, ack => convTranspose_CP_34_elements(90)); -- 
    cr_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(90), ack => RPIPE_ConvTranspose_input_pipe_300_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_300_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Sample/rr
      -- 
    ca_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_300_inst_ack_1, ack => convTranspose_CP_34_elements(91)); -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => type_cast_304_inst_req_0); -- 
    rr_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => RPIPE_ConvTranspose_input_pipe_312_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Sample/ra
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_304_inst_ack_0, ack => convTranspose_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_304_Update/ca
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_304_inst_ack_1, ack => convTranspose_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_update_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Update/cr
      -- 
    ra_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_312_inst_ack_0, ack => convTranspose_CP_34_elements(94)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(94), ack => RPIPE_ConvTranspose_input_pipe_312_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_312_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Sample/rr
      -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_312_inst_ack_1, ack => convTranspose_CP_34_elements(95)); -- 
    rr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => type_cast_316_inst_req_0); -- 
    rr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => RPIPE_ConvTranspose_input_pipe_325_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Sample/ra
      -- 
    ra_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_0, ack => convTranspose_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_316_Update/ca
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_1, ack => convTranspose_CP_34_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_update_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Update/cr
      -- 
    ra_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_325_inst_ack_0, ack => convTranspose_CP_34_elements(98)); -- 
    cr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(98), ack => RPIPE_ConvTranspose_input_pipe_325_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_325_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Sample/rr
      -- 
    ca_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_325_inst_ack_1, ack => convTranspose_CP_34_elements(99)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => type_cast_329_inst_req_0); -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => RPIPE_ConvTranspose_input_pipe_337_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Sample/ra
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_329_inst_ack_0, ack => convTranspose_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_329_Update/ca
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_329_inst_ack_1, ack => convTranspose_CP_34_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_update_start_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Update/cr
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_337_inst_ack_0, ack => convTranspose_CP_34_elements(102)); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(102), ack => RPIPE_ConvTranspose_input_pipe_337_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_337_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Sample/rr
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_337_inst_ack_1, ack => convTranspose_CP_34_elements(103)); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => type_cast_341_inst_req_0); -- 
    rr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => RPIPE_ConvTranspose_input_pipe_350_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Sample/ra
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_341_inst_ack_0, ack => convTranspose_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_341_Update/ca
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_341_inst_ack_1, ack => convTranspose_CP_34_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_update_start_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Update/cr
      -- 
    ra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_350_inst_ack_0, ack => convTranspose_CP_34_elements(106)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(106), ack => RPIPE_ConvTranspose_input_pipe_350_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_350_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Sample/rr
      -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_350_inst_ack_1, ack => convTranspose_CP_34_elements(107)); -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => type_cast_354_inst_req_0); -- 
    rr_846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => RPIPE_ConvTranspose_input_pipe_362_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Sample/ra
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_354_inst_ack_0, ack => convTranspose_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_354_Update/ca
      -- 
    ca_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_354_inst_ack_1, ack => convTranspose_CP_34_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_update_start_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Update/cr
      -- 
    ra_847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_362_inst_ack_0, ack => convTranspose_CP_34_elements(110)); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(110), ack => RPIPE_ConvTranspose_input_pipe_362_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_362_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Sample/rr
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_362_inst_ack_1, ack => convTranspose_CP_34_elements(111)); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => RPIPE_ConvTranspose_input_pipe_375_inst_req_0); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => type_cast_366_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Sample/ra
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_366_inst_ack_0, ack => convTranspose_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_366_Update/ca
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_366_inst_ack_1, ack => convTranspose_CP_34_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_update_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Update/cr
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_375_inst_ack_0, ack => convTranspose_CP_34_elements(114)); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(114), ack => RPIPE_ConvTranspose_input_pipe_375_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/RPIPE_ConvTranspose_input_pipe_375_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Sample/rr
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_375_inst_ack_1, ack => convTranspose_CP_34_elements(115)); -- 
    rr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(115), ack => type_cast_379_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Sample/ra
      -- 
    ra_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_379_inst_ack_0, ack => convTranspose_CP_34_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/type_cast_379_Update/ca
      -- 
    ca_894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_379_inst_ack_1, ack => convTranspose_CP_34_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391__exit__
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392__entry__
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_391/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_32/R_cmp456_393_place
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_392_else_link/$entry
      -- 
    branch_req_902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(118), ack => if_stmt_392_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(117) & convTranspose_CP_34_elements(105) & convTranspose_CP_34_elements(113) & convTranspose_CP_34_elements(89) & convTranspose_CP_34_elements(109) & convTranspose_CP_34_elements(93) & convTranspose_CP_34_elements(97) & convTranspose_CP_34_elements(101) & convTranspose_CP_34_elements(85) & convTranspose_CP_34_elements(59) & convTranspose_CP_34_elements(62) & convTranspose_CP_34_elements(65) & convTranspose_CP_34_elements(68) & convTranspose_CP_34_elements(71) & convTranspose_CP_34_elements(74) & convTranspose_CP_34_elements(77) & convTranspose_CP_34_elements(81);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_413__exit__
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448__entry__
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_392_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_392_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph458
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_update_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph458_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph458_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_413_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_413_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_413_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_413_PhiAck/dummy
      -- 
    if_choice_transition_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_392_branch_ack_1, ack => convTranspose_CP_34_elements(119)); -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_434_inst_req_0); -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_434_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	360 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_392_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_392_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_392_branch_ack_0, ack => convTranspose_CP_34_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	360 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_620__exit__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655__entry__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_update_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_407_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_407_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph454
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph454_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph454_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_620_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_620_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_620_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_620_PhiAck/dummy
      -- 
    if_choice_transition_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_407_branch_ack_1, ack => convTranspose_CP_34_elements(121)); -- 
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_641_inst_req_1); -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_641_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	360 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	373 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_407_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_407_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_407_branch_ack_0, ack => convTranspose_CP_34_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Sample/ra
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_434_inst_ack_0, ack => convTranspose_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	361 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448__exit__
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_419_to_assign_stmt_448/type_cast_434_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_451/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/$entry
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_434_inst_ack_1, ack => convTranspose_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	366 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_sample_complete
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_463_index_offset_ack_0, ack => convTranspose_CP_34_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	366 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_request/req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Update/$exit
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_463_index_offset_ack_1, ack => convTranspose_CP_34_elements(126)); -- 
    req_995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(126), ack => addr_of_464_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_request/ack
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_request/$exit
      -- 
    ack_996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_464_final_reg_ack_0, ack => convTranspose_CP_34_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	366 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_complete/ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_complete/$exit
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_464_final_reg_ack_1, ack => convTranspose_CP_34_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	366 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_update_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_sample_completed_
      -- 
    ra_1010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_467_inst_ack_0, ack => convTranspose_CP_34_elements(129)); -- 
    cr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(129), ack => RPIPE_ConvTranspose_input_pipe_467_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_update_completed_
      -- 
    ca_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_467_inst_ack_1, ack => convTranspose_CP_34_elements(130)); -- 
    rr_1023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => type_cast_471_inst_req_0); -- 
    rr_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => RPIPE_ConvTranspose_input_pipe_480_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_sample_completed_
      -- 
    ra_1024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_471_inst_ack_0, ack => convTranspose_CP_34_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	366 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_update_completed_
      -- 
    ca_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_471_inst_ack_1, ack => convTranspose_CP_34_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_update_start_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_sample_completed_
      -- 
    ra_1038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_480_inst_ack_0, ack => convTranspose_CP_34_elements(133)); -- 
    cr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(133), ack => RPIPE_ConvTranspose_input_pipe_480_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_480_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Sample/$entry
      -- 
    ca_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_480_inst_ack_1, ack => convTranspose_CP_34_elements(134)); -- 
    rr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => type_cast_484_inst_req_0); -- 
    rr_1065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_sample_completed_
      -- 
    ra_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_484_inst_ack_0, ack => convTranspose_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	366 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_update_completed_
      -- 
    ca_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_484_inst_ack_1, ack => convTranspose_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_update_start_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_sample_completed_
      -- 
    ra_1066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_0, ack => convTranspose_CP_34_elements(137)); -- 
    cr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(137), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_498_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Sample/$entry
      -- 
    ca_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_1, ack => convTranspose_CP_34_elements(138)); -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => type_cast_502_inst_req_0); -- 
    rr_1093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_sample_completed_
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_0, ack => convTranspose_CP_34_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	366 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_update_completed_
      -- 
    ca_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_1, ack => convTranspose_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_update_start_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_sample_completed_
      -- 
    ra_1094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_0, ack => convTranspose_CP_34_elements(141)); -- 
    cr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(141), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_516_update_completed_
      -- 
    ca_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_1, ack => convTranspose_CP_34_elements(142)); -- 
    rr_1107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => type_cast_520_inst_req_0); -- 
    rr_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_sample_completed_
      -- 
    ra_1108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => convTranspose_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	366 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_update_completed_
      -- 
    ca_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => convTranspose_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_update_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_sample_completed_
      -- 
    ra_1122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_0, ack => convTranspose_CP_34_elements(145)); -- 
    cr_1126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(145), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_534_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_sample_start_
      -- 
    ca_1127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_1, ack => convTranspose_CP_34_elements(146)); -- 
    rr_1135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => type_cast_538_inst_req_0); -- 
    rr_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Sample/ra
      -- 
    ra_1136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convTranspose_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	366 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Update/$exit
      -- 
    ca_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convTranspose_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_update_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_sample_completed_
      -- 
    ra_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_0, ack => convTranspose_CP_34_elements(149)); -- 
    cr_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(149), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_552_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Sample/$entry
      -- 
    ca_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_1, ack => convTranspose_CP_34_elements(150)); -- 
    rr_1163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => type_cast_556_inst_req_0); -- 
    rr_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_sample_completed_
      -- 
    ra_1164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_0, ack => convTranspose_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	366 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_update_completed_
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_1, ack => convTranspose_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_update_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Sample/$exit
      -- 
    ra_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_0, ack => convTranspose_CP_34_elements(153)); -- 
    cr_1182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(153), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_570_update_completed_
      -- 
    ca_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_1, ack => convTranspose_CP_34_elements(154)); -- 
    rr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => type_cast_574_inst_req_0); -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_sample_completed_
      -- 
    ra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_0, ack => convTranspose_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	366 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_update_completed_
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_1, ack => convTranspose_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_update_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Update/$entry
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_0, ack => convTranspose_CP_34_elements(157)); -- 
    cr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(157), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_588_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Sample/$entry
      -- 
    ca_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_1, ack => convTranspose_CP_34_elements(158)); -- 
    rr_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(158), ack => type_cast_592_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Sample/ra
      -- 
    ra_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => convTranspose_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	366 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_update_completed_
      -- 
    ca_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => convTranspose_CP_34_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/ptr_deref_600_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/ptr_deref_600_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/ptr_deref_600_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/ptr_deref_600_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/$entry
      -- 
    rr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(161), ack => ptr_deref_600_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(128) & convTranspose_CP_34_elements(132) & convTranspose_CP_34_elements(136) & convTranspose_CP_34_elements(140) & convTranspose_CP_34_elements(144) & convTranspose_CP_34_elements(148) & convTranspose_CP_34_elements(152) & convTranspose_CP_34_elements(156) & convTranspose_CP_34_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Sample/$exit
      -- 
    ra_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_store_0_ack_0, ack => convTranspose_CP_34_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	366 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/word_access_complete/word_0/$exit
      -- 
    ca_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_store_0_ack_1, ack => convTranspose_CP_34_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	125 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613__exit__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614__entry__
      -- CP-element group 164: 	 branch_block_stmt_32/R_exitcond3_615_place
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_614_else_link/$entry
      -- 
    branch_req_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(164), ack => if_stmt_614_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(125) & convTranspose_CP_34_elements(163);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	360 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_614_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_398__exit__
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_614_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_398_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_398_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_398_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_398_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_614_branch_ack_1, ack => convTranspose_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	362 
    -- CP-element group 166: 	363 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_614_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_614_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_614_branch_ack_0, ack => convTranspose_CP_34_elements(166)); -- 
    rr_2797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_457_inst_req_0); -- 
    cr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_457_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_sample_completed_
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_0, ack => convTranspose_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	367 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655__exit__
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_626_to_assign_stmt_655/type_cast_641_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_658/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/$entry
      -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_1, ack => convTranspose_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	372 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_sample_complete
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_670_index_offset_ack_0, ack => convTranspose_CP_34_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	372 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_request/req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Update/$exit
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_670_index_offset_ack_1, ack => convTranspose_CP_34_elements(170)); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(170), ack => addr_of_671_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_request/ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_sample_completed_
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_671_final_reg_ack_0, ack => convTranspose_CP_34_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	372 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_word_addrgen/root_register_ack
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_671_final_reg_ack_1, ack => convTranspose_CP_34_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	372 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_update_start_
      -- 
    ra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_674_inst_ack_0, ack => convTranspose_CP_34_elements(173)); -- 
    cr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(173), ack => RPIPE_ConvTranspose_input_pipe_674_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Sample/$entry
      -- 
    ca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_674_inst_ack_1, ack => convTranspose_CP_34_elements(174)); -- 
    rr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => type_cast_678_inst_req_0); -- 
    rr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => RPIPE_ConvTranspose_input_pipe_687_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Sample/$exit
      -- 
    ra_1383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_678_inst_ack_0, ack => convTranspose_CP_34_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	372 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Update/$exit
      -- 
    ca_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_678_inst_ack_1, ack => convTranspose_CP_34_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_update_start_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_sample_completed_
      -- 
    ra_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_687_inst_ack_0, ack => convTranspose_CP_34_elements(177)); -- 
    cr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(177), ack => RPIPE_ConvTranspose_input_pipe_687_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_687_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Sample/rr
      -- 
    ca_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_687_inst_ack_1, ack => convTranspose_CP_34_elements(178)); -- 
    rr_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => type_cast_691_inst_req_0); -- 
    rr_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_sample_completed_
      -- 
    ra_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_0, ack => convTranspose_CP_34_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	372 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_update_completed_
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_1, ack => convTranspose_CP_34_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_update_start_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Update/cr
      -- 
    ra_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_0, ack => convTranspose_CP_34_elements(181)); -- 
    cr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(181), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_705_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Sample/rr
      -- 
    ca_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_1, ack => convTranspose_CP_34_elements(182)); -- 
    rr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => type_cast_709_inst_req_0); -- 
    rr_1452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Sample/ra
      -- 
    ra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => convTranspose_CP_34_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	372 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Update/ca
      -- 
    ca_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => convTranspose_CP_34_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_update_start_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Update/cr
      -- 
    ra_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_0, ack => convTranspose_CP_34_elements(185)); -- 
    cr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(185), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_723_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Sample/rr
      -- 
    ca_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_1, ack => convTranspose_CP_34_elements(186)); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => type_cast_727_inst_req_0); -- 
    rr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Sample/ra
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => convTranspose_CP_34_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	372 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Update/ca
      -- 
    ca_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => convTranspose_CP_34_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_update_start_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Update/cr
      -- 
    ra_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_0, ack => convTranspose_CP_34_elements(189)); -- 
    cr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(189), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_741_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Sample/rr
      -- 
    ca_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_1, ack => convTranspose_CP_34_elements(190)); -- 
    rr_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => type_cast_745_inst_req_0); -- 
    rr_1508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Sample/ra
      -- 
    ra_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_0, ack => convTranspose_CP_34_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	372 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Update/ca
      -- 
    ca_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_1, ack => convTranspose_CP_34_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_update_start_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Update/cr
      -- 
    ra_1509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_0, ack => convTranspose_CP_34_elements(193)); -- 
    cr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(193), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_759_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Sample/rr
      -- 
    ca_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_1, ack => convTranspose_CP_34_elements(194)); -- 
    rr_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => type_cast_763_inst_req_0); -- 
    rr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Sample/ra
      -- 
    ra_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => convTranspose_CP_34_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	372 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Update/ca
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_1, ack => convTranspose_CP_34_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_update_start_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Update/cr
      -- 
    ra_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_0, ack => convTranspose_CP_34_elements(197)); -- 
    cr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(197), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_777_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Sample/rr
      -- 
    ca_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_1, ack => convTranspose_CP_34_elements(198)); -- 
    rr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => type_cast_781_inst_req_0); -- 
    rr_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Sample/ra
      -- 
    ra_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => convTranspose_CP_34_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	372 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Update/ca
      -- 
    ca_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => convTranspose_CP_34_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_update_start_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Update/cr
      -- 
    ra_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_0, ack => convTranspose_CP_34_elements(201)); -- 
    cr_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(201), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_795_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Sample/rr
      -- 
    ca_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_1, ack => convTranspose_CP_34_elements(202)); -- 
    rr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(202), ack => type_cast_799_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Sample/ra
      -- 
    ra_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => convTranspose_CP_34_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	372 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Update/ca
      -- 
    ca_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => convTranspose_CP_34_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/ptr_deref_807_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/ptr_deref_807_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/ptr_deref_807_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/ptr_deref_807_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/word_access_start/word_0/rr
      -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(205), ack => ptr_deref_807_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(204) & convTranspose_CP_34_elements(172) & convTranspose_CP_34_elements(176) & convTranspose_CP_34_elements(180) & convTranspose_CP_34_elements(184) & convTranspose_CP_34_elements(188) & convTranspose_CP_34_elements(192) & convTranspose_CP_34_elements(196) & convTranspose_CP_34_elements(200);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Sample/word_access_start/word_0/ra
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_store_0_ack_0, ack => convTranspose_CP_34_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	372 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/word_access_complete/word_0/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_store_0_ack_1, ack => convTranspose_CP_34_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820__exit__
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821__entry__
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_32/R_exitcond2_822_place
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_821_else_link/$entry
      -- 
    branch_req_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(208), ack => if_stmt_821_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(207) & convTranspose_CP_34_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	373 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_827__exit__
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_821_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_821_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_827_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_827_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_827_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_827_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_821_branch_ack_1, ack => convTranspose_CP_34_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	368 
    -- CP-element group 210: 	369 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_821_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_821_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_821_branch_ack_0, ack => convTranspose_CP_34_elements(210)); -- 
    rr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_664_inst_req_0); -- 
    cr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_664_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	373 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Sample/ra
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_0, ack => convTranspose_CP_34_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	373 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Update/ca
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_1, ack => convTranspose_CP_34_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	373 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_836_inst_ack_0, ack => convTranspose_CP_34_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	373 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_836_inst_ack_1, ack => convTranspose_CP_34_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	373 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_840_inst_ack_0, ack => convTranspose_CP_34_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	373 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_840_inst_ack_1, ack => convTranspose_CP_34_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857__exit__
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858__entry__
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_32/R_cmp264448_859_place
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_858_else_link/$entry
      -- 
    branch_req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(217), ack => if_stmt_858_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(212) & convTranspose_CP_34_elements(214) & convTranspose_CP_34_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_864__exit__
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899__entry__
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_858_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_858_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph450
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_update_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph450_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph450_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_864_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_864_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_864_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_864_PhiAck/dummy
      -- 
    if_choice_transition_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_858_branch_ack_1, ack => convTranspose_CP_34_elements(218)); -- 
    rr_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_885_inst_req_0); -- 
    cr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_885_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	380 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_858_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_858_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273
      -- 
    else_choice_transition_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_858_branch_ack_0, ack => convTranspose_CP_34_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Sample/ra
      -- 
    ra_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_885_inst_ack_0, ack => convTranspose_CP_34_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	374 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_870_to_assign_stmt_899/type_cast_885_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_902/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/$entry
      -- 
    ca_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_885_inst_ack_1, ack => convTranspose_CP_34_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	379 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Sample/ack
      -- 
    ack_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_offset_ack_0, ack => convTranspose_CP_34_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	379 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_request/req
      -- 
    ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_offset_ack_1, ack => convTranspose_CP_34_elements(223)); -- 
    req_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(223), ack => addr_of_915_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_request/ack
      -- 
    ack_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_915_final_reg_ack_0, ack => convTranspose_CP_34_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	379 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/ptr_deref_918_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/ptr_deref_918_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/ptr_deref_918_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/ptr_deref_918_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/word_access_start/word_0/rr
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_915_final_reg_ack_1, ack => convTranspose_CP_34_elements(225)); -- 
    rr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(225), ack => ptr_deref_918_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Sample/word_access_start/word_0/ra
      -- 
    ra_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_918_store_0_ack_0, ack => convTranspose_CP_34_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	379 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/word_access_complete/word_0/ca
      -- 
    ca_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_918_store_0_ack_1, ack => convTranspose_CP_34_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: 	222 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932__exit__
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933__entry__
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_32/R_exitcond_934_place
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_933_else_link/$entry
      -- 
    branch_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(228), ack => if_stmt_933_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(227) & convTranspose_CP_34_elements(222);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	380 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_939__exit__
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_939_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_939_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_939_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_939_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_933_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_933_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit
      -- 
    if_choice_transition_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_933_branch_ack_1, ack => convTranspose_CP_34_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	375 
    -- CP-element group 230: 	376 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Update/cr
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_933_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_933_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- 
    else_choice_transition_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_933_branch_ack_0, ack => convTranspose_CP_34_elements(230)); -- 
    rr_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_908_inst_req_0); -- 
    cr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_908_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	380 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Sample/cra
      -- 
    cra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_944_call_ack_0, ack => convTranspose_CP_34_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	380 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Sample/rr
      -- 
    cca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_944_call_ack_1, ack => convTranspose_CP_34_elements(232)); -- 
    rr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(232), ack => type_cast_949_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Sample/ra
      -- 
    ra_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_949_inst_ack_0, ack => convTranspose_CP_34_elements(233)); -- 
    -- CP-element group 234:  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	380 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (10) 
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950__exit__
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995__entry__
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Sample/req
      -- 
    ca_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_949_inst_ack_1, ack => convTranspose_CP_34_elements(234)); -- 
    req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block0_start_952_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_update_start_
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Update/req
      -- 
    ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_952_inst_ack_0, ack => convTranspose_CP_34_elements(235)); -- 
    req_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(235), ack => WPIPE_Block0_start_952_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_952_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Sample/req
      -- 
    ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_952_inst_ack_1, ack => convTranspose_CP_34_elements(236)); -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(236), ack => WPIPE_Block0_start_955_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Update/req
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_955_inst_ack_0, ack => convTranspose_CP_34_elements(237)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(237), ack => WPIPE_Block0_start_955_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_955_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Sample/req
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_955_inst_ack_1, ack => convTranspose_CP_34_elements(238)); -- 
    req_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(238), ack => WPIPE_Block0_start_958_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_update_start_
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Update/req
      -- 
    ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_958_inst_ack_0, ack => convTranspose_CP_34_elements(239)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(239), ack => WPIPE_Block0_start_958_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_958_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Sample/req
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_958_inst_ack_1, ack => convTranspose_CP_34_elements(240)); -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(240), ack => WPIPE_Block0_start_961_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Update/req
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_961_inst_ack_0, ack => convTranspose_CP_34_elements(241)); -- 
    req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(241), ack => WPIPE_Block0_start_961_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_961_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Sample/req
      -- 
    ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_961_inst_ack_1, ack => convTranspose_CP_34_elements(242)); -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(242), ack => WPIPE_Block0_start_964_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_update_start_
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Update/req
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_964_inst_ack_0, ack => convTranspose_CP_34_elements(243)); -- 
    req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(243), ack => WPIPE_Block0_start_964_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_964_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Sample/req
      -- 
    ack_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_964_inst_ack_1, ack => convTranspose_CP_34_elements(244)); -- 
    req_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(244), ack => WPIPE_Block0_start_967_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_update_start_
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Update/req
      -- 
    ack_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_967_inst_ack_0, ack => convTranspose_CP_34_elements(245)); -- 
    req_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(245), ack => WPIPE_Block0_start_967_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_967_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Sample/req
      -- 
    ack_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_967_inst_ack_1, ack => convTranspose_CP_34_elements(246)); -- 
    req_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(246), ack => WPIPE_Block0_start_970_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Update/req
      -- 
    ack_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_0, ack => convTranspose_CP_34_elements(247)); -- 
    req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(247), ack => WPIPE_Block0_start_970_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_970_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Sample/req
      -- 
    ack_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_1, ack => convTranspose_CP_34_elements(248)); -- 
    req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(248), ack => WPIPE_Block0_start_973_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Update/req
      -- 
    ack_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_0, ack => convTranspose_CP_34_elements(249)); -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(249), ack => WPIPE_Block0_start_973_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_973_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Sample/req
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_1, ack => convTranspose_CP_34_elements(250)); -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(250), ack => WPIPE_Block0_start_976_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_update_start_
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Update/req
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_0, ack => convTranspose_CP_34_elements(251)); -- 
    req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(251), ack => WPIPE_Block0_start_976_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_976_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Sample/req
      -- 
    ack_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_1, ack => convTranspose_CP_34_elements(252)); -- 
    req_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(252), ack => WPIPE_Block0_start_979_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Update/req
      -- 
    ack_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_0, ack => convTranspose_CP_34_elements(253)); -- 
    req_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(253), ack => WPIPE_Block0_start_979_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_979_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Sample/req
      -- 
    ack_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_1, ack => convTranspose_CP_34_elements(254)); -- 
    req_2034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(254), ack => WPIPE_Block0_start_983_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Sample/ack
      -- 
    ack_2035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_0, ack => convTranspose_CP_34_elements(255)); -- 
    req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(255), ack => WPIPE_Block0_start_983_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_983_update_completed_
      -- 
    ack_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_1, ack => convTranspose_CP_34_elements(256)); -- 
    req_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(256), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_update_start_
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Update/req
      -- 
    ack_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_34_elements(257)); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(257), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_987_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Sample/req
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_34_elements(258)); -- 
    req_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(258), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Sample/$exit
      -- 
    ack_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_34_elements(259)); -- 
    req_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(259), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_990_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Sample/req
      -- 
    ack_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_34_elements(260)); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(260), ack => WPIPE_Block0_start_993_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Update/req
      -- 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_0, ack => convTranspose_CP_34_elements(261)); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(261), ack => WPIPE_Block0_start_993_inst_req_1); -- 
    -- CP-element group 262:  transition  place  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (10) 
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995__exit__
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_999__entry__
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_999/$entry
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/WPIPE_Block0_start_993_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_954_to_assign_stmt_995/$exit
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_1, ack => convTranspose_CP_34_elements(262)); -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(262), ack => RPIPE_Block0_done_998_inst_req_0); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Sample/ra
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_update_start_
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_sample_completed_
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_998_inst_ack_0, ack => convTranspose_CP_34_elements(263)); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(263), ack => RPIPE_Block0_done_998_inst_req_1); -- 
    -- CP-element group 264:  fork  transition  place  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264: 	266 
    -- CP-element group 264: 	268 
    -- CP-element group 264: 	270 
    -- CP-element group 264: 	272 
    -- CP-element group 264: 	274 
    -- CP-element group 264: 	276 
    -- CP-element group 264: 	278 
    -- CP-element group 264: 	280 
    -- CP-element group 264: 	282 
    -- CP-element group 264: 	284 
    -- CP-element group 264:  members (40) 
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_999__exit__
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110__entry__
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Update/ccr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Sample/crr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Update/ca
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_999/RPIPE_Block0_done_998_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_999/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_update_start_
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_998_inst_ack_1, ack => convTranspose_CP_34_elements(264)); -- 
    cr_2143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1015_inst_req_1); -- 
    ccr_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => call_stmt_1002_call_req_1); -- 
    crr_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => call_stmt_1002_call_req_0); -- 
    cr_2213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1065_inst_req_1); -- 
    cr_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1055_inst_req_1); -- 
    cr_2227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1075_inst_req_1); -- 
    cr_2129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1006_inst_req_1); -- 
    cr_2185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1045_inst_req_1); -- 
    cr_2171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1035_inst_req_1); -- 
    cr_2241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1085_inst_req_1); -- 
    cr_2157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => type_cast_1025_inst_req_1); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Sample/cra
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_sample_completed_
      -- 
    cra_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1002_call_ack_0, ack => convTranspose_CP_34_elements(265)); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_Update/cca
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Sample/rr
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/call_stmt_1002_update_completed_
      -- 
    cca_2116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1002_call_ack_1, ack => convTranspose_CP_34_elements(266)); -- 
    rr_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(266), ack => type_cast_1006_inst_req_0); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Sample/ra
      -- 
    ra_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1006_inst_ack_0, ack => convTranspose_CP_34_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	264 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	271 
    -- CP-element group 268: 	273 
    -- CP-element group 268: 	275 
    -- CP-element group 268: 	277 
    -- CP-element group 268: 	279 
    -- CP-element group 268: 	281 
    -- CP-element group 268: 	283 
    -- CP-element group 268:  members (27) 
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1006_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Sample/$entry
      -- 
    ca_2130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1006_inst_ack_1, ack => convTranspose_CP_34_elements(268)); -- 
    rr_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1015_inst_req_0); -- 
    rr_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1025_inst_req_0); -- 
    rr_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1035_inst_req_0); -- 
    rr_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1045_inst_req_0); -- 
    rr_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1055_inst_req_0); -- 
    rr_2208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1065_inst_req_0); -- 
    rr_2222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1075_inst_req_0); -- 
    rr_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => type_cast_1085_inst_req_0); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Sample/ra
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_sample_completed_
      -- 
    ra_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_0, ack => convTranspose_CP_34_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	264 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	305 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Update/ca
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1015_update_completed_
      -- 
    ca_2144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_1, ack => convTranspose_CP_34_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	268 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Sample/ra
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Sample/$exit
      -- 
    ra_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_0, ack => convTranspose_CP_34_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	264 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	302 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Update/ca
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1025_update_completed_
      -- 
    ca_2158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_1, ack => convTranspose_CP_34_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	268 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Sample/ra
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_sample_completed_
      -- 
    ra_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_0, ack => convTranspose_CP_34_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	264 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	299 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Update/ca
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1035_update_completed_
      -- 
    ca_2172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_1, ack => convTranspose_CP_34_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	268 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_sample_completed_
      -- 
    ra_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_0, ack => convTranspose_CP_34_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	264 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	296 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1045_update_completed_
      -- 
    ca_2186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_1, ack => convTranspose_CP_34_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	268 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Sample/ra
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_sample_completed_
      -- 
    ra_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => convTranspose_CP_34_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	264 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	293 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1055_update_completed_
      -- 
    ca_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => convTranspose_CP_34_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	268 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Sample/$exit
      -- 
    ra_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_0, ack => convTranspose_CP_34_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	264 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	290 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_Update/ca
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1065_update_completed_
      -- 
    ca_2214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_1, ack => convTranspose_CP_34_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	268 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Sample/$exit
      -- 
    ra_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1075_inst_ack_0, ack => convTranspose_CP_34_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	264 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	287 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1075_Update/ca
      -- 
    ca_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1075_inst_ack_1, ack => convTranspose_CP_34_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	268 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Sample/ra
      -- 
    ra_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_0, ack => convTranspose_CP_34_elements(283)); -- 
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	264 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Sample/req
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Update/ca
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/type_cast_1085_Update/$exit
      -- 
    ca_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_1, ack => convTranspose_CP_34_elements(284)); -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(284), ack => WPIPE_ConvTranspose_output_pipe_1087_inst_req_0); -- 
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Update/req
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_update_start_
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_sample_completed_
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1087_inst_ack_0, ack => convTranspose_CP_34_elements(285)); -- 
    req_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(285), ack => WPIPE_ConvTranspose_output_pipe_1087_inst_req_1); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1087_update_completed_
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1087_inst_ack_1, ack => convTranspose_CP_34_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	282 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Sample/req
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Sample/$entry
      -- 
    req_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(287), ack => WPIPE_ConvTranspose_output_pipe_1090_inst_req_0); -- 
    convTranspose_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(282) & convTranspose_CP_34_elements(286);
      gj_convTranspose_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_update_start_
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Sample/ack
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Update/req
      -- 
    ack_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1090_inst_ack_0, ack => convTranspose_CP_34_elements(288)); -- 
    req_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(288), ack => WPIPE_ConvTranspose_output_pipe_1090_inst_req_1); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1090_Update/ack
      -- 
    ack_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1090_inst_ack_1, ack => convTranspose_CP_34_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	280 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_sample_start_
      -- 
    req_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(290), ack => WPIPE_ConvTranspose_output_pipe_1093_inst_req_0); -- 
    convTranspose_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(280) & convTranspose_CP_34_elements(289);
      gj_convTranspose_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Update/req
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_update_start_
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_sample_completed_
      -- 
    ack_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1093_inst_ack_0, ack => convTranspose_CP_34_elements(291)); -- 
    req_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(291), ack => WPIPE_ConvTranspose_output_pipe_1093_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1093_update_completed_
      -- 
    ack_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1093_inst_ack_1, ack => convTranspose_CP_34_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	278 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_sample_start_
      -- 
    req_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(293), ack => WPIPE_ConvTranspose_output_pipe_1096_inst_req_0); -- 
    convTranspose_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(278) & convTranspose_CP_34_elements(292);
      gj_convTranspose_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Update/req
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_update_start_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_sample_completed_
      -- 
    ack_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1096_inst_ack_0, ack => convTranspose_CP_34_elements(294)); -- 
    req_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(294), ack => WPIPE_ConvTranspose_output_pipe_1096_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_Update/ack
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1096_update_completed_
      -- 
    ack_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1096_inst_ack_1, ack => convTranspose_CP_34_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	276 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Sample/req
      -- 
    req_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(296), ack => WPIPE_ConvTranspose_output_pipe_1099_inst_req_0); -- 
    convTranspose_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(276) & convTranspose_CP_34_elements(295);
      gj_convTranspose_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_update_start_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Update/req
      -- 
    ack_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1099_inst_ack_0, ack => convTranspose_CP_34_elements(297)); -- 
    req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(297), ack => WPIPE_ConvTranspose_output_pipe_1099_inst_req_1); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1099_Update/ack
      -- 
    ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1099_inst_ack_1, ack => convTranspose_CP_34_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	274 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Sample/req
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_sample_start_
      -- 
    req_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(299), ack => WPIPE_ConvTranspose_output_pipe_1102_inst_req_0); -- 
    convTranspose_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(274) & convTranspose_CP_34_elements(298);
      gj_convTranspose_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Update/req
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Sample/ack
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_update_start_
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_sample_completed_
      -- 
    ack_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1102_inst_ack_0, ack => convTranspose_CP_34_elements(300)); -- 
    req_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(300), ack => WPIPE_ConvTranspose_output_pipe_1102_inst_req_1); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_Update/ack
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1102_update_completed_
      -- 
    ack_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1102_inst_ack_1, ack => convTranspose_CP_34_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	272 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Sample/$entry
      -- 
    req_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(302), ack => WPIPE_ConvTranspose_output_pipe_1105_inst_req_0); -- 
    convTranspose_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(272) & convTranspose_CP_34_elements(301);
      gj_convTranspose_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Update/req
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Sample/$exit
      -- 
    ack_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1105_inst_ack_0, ack => convTranspose_CP_34_elements(303)); -- 
    req_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(303), ack => WPIPE_ConvTranspose_output_pipe_1105_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1105_Update/$exit
      -- 
    ack_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1105_inst_ack_1, ack => convTranspose_CP_34_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	270 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Sample/req
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Sample/$entry
      -- 
    req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(305), ack => WPIPE_ConvTranspose_output_pipe_1108_inst_req_0); -- 
    convTranspose_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(270) & convTranspose_CP_34_elements(304);
      gj_convTranspose_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_update_start_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Update/req
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Sample/ack
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Sample/$exit
      -- 
    ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1108_inst_ack_0, ack => convTranspose_CP_34_elements(306)); -- 
    req_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(306), ack => WPIPE_ConvTranspose_output_pipe_1108_inst_req_1); -- 
    -- CP-element group 307:  branch  transition  place  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (13) 
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112_dead_link/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110__exit__
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112__entry__
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/WPIPE_ConvTranspose_output_pipe_1108_Update/ack
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112_eval_test/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112_else_link/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_1002_to_assign_stmt_1110/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112_if_link/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/R_cmp264448_1113_place
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112_eval_test/branch_req
      -- CP-element group 307: 	 branch_block_stmt_32/if_stmt_1112_eval_test/$exit
      -- 
    ack_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1108_inst_ack_1, ack => convTranspose_CP_34_elements(307)); -- 
    branch_req_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(307), ack => if_stmt_1112_branch_req_0); -- 
    -- CP-element group 308:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	310 
    -- CP-element group 308: 	311 
    -- CP-element group 308:  members (18) 
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1118__exit__
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153__entry__
      -- CP-element group 308: 	 branch_block_stmt_32/forx_xend273_bbx_xnph
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1118_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Sample/rr
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_update_start_
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_32/if_stmt_1112_if_link/if_choice_transition
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/if_stmt_1112_if_link/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1118_PhiAck/dummy
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1118_PhiAck/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1118_PhiAck/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$entry
      -- 
    if_choice_transition_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1112_branch_ack_1, ack => convTranspose_CP_34_elements(308)); -- 
    rr_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(308), ack => type_cast_1139_inst_req_0); -- 
    cr_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(308), ack => type_cast_1139_inst_req_1); -- 
    -- CP-element group 309:  transition  place  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	387 
    -- CP-element group 309:  members (5) 
      -- CP-element group 309: 	 branch_block_stmt_32/forx_xend273_forx_xend443_PhiReq/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/if_stmt_1112_else_link/else_choice_transition
      -- CP-element group 309: 	 branch_block_stmt_32/forx_xend273_forx_xend443
      -- CP-element group 309: 	 branch_block_stmt_32/if_stmt_1112_else_link/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/forx_xend273_forx_xend443_PhiReq/$entry
      -- 
    else_choice_transition_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1112_branch_ack_0, ack => convTranspose_CP_34_elements(309)); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Sample/ra
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_sample_completed_
      -- 
    ra_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1139_inst_ack_0, ack => convTranspose_CP_34_elements(310)); -- 
    -- CP-element group 311:  transition  place  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	308 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	381 
    -- CP-element group 311:  members (9) 
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153__exit__
      -- CP-element group 311: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Update/ca
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/type_cast_1139_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_1124_to_assign_stmt_1153/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1156/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/$entry
      -- 
    ca_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1139_inst_ack_1, ack => convTranspose_CP_34_elements(311)); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	386 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	357 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_sample_complete
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Sample/ack
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1168_index_offset_ack_0, ack => convTranspose_CP_34_elements(312)); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	386 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (11) 
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_offset_calculated
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_root_address_calculated
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_base_plus_offset/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_base_plus_offset/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_base_plus_offset/sum_rename_req
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_base_plus_offset/sum_rename_ack
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_request/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_request/req
      -- 
    ack_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1168_index_offset_ack_1, ack => convTranspose_CP_34_elements(313)); -- 
    req_2433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(313), ack => addr_of_1169_final_reg_req_0); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_request/$exit
      -- CP-element group 314: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_request/ack
      -- 
    ack_2434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1169_final_reg_ack_0, ack => convTranspose_CP_34_elements(314)); -- 
    -- CP-element group 315:  join  fork  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	386 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (24) 
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_complete/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_complete/ack
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_sample_start_
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_address_calculated
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_word_address_calculated
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_root_address_calculated
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_address_resized
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_addr_resize/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_addr_resize/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_addr_resize/base_resize_req
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_addr_resize/base_resize_ack
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_plus_offset/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_plus_offset/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_plus_offset/sum_rename_req
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_base_plus_offset/sum_rename_ack
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_word_addrgen/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_word_addrgen/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_word_addrgen/root_register_req
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_word_addrgen/root_register_ack
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/word_access_start/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/word_access_start/word_0/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/word_access_start/word_0/rr
      -- 
    ack_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1169_final_reg_ack_1, ack => convTranspose_CP_34_elements(315)); -- 
    rr_2472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(315), ack => ptr_deref_1173_load_0_req_0); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (5) 
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_sample_completed_
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/word_access_start/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/word_access_start/word_0/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Sample/word_access_start/word_0/ra
      -- 
    ra_2473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1173_load_0_ack_0, ack => convTranspose_CP_34_elements(316)); -- 
    -- CP-element group 317:  fork  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	386 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317: 	320 
    -- CP-element group 317: 	322 
    -- CP-element group 317: 	324 
    -- CP-element group 317: 	326 
    -- CP-element group 317: 	328 
    -- CP-element group 317: 	330 
    -- CP-element group 317: 	332 
    -- CP-element group 317:  members (33) 
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/word_access_complete/$exit
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/word_access_complete/word_0/$exit
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/word_access_complete/word_0/ca
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/ptr_deref_1173_Merge/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/ptr_deref_1173_Merge/$exit
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/ptr_deref_1173_Merge/merge_req
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/ptr_deref_1173_Merge/merge_ack
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Sample/rr
      -- 
    ca_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1173_load_0_ack_1, ack => convTranspose_CP_34_elements(317)); -- 
    rr_2497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1177_inst_req_0); -- 
    rr_2511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1187_inst_req_0); -- 
    rr_2525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1197_inst_req_0); -- 
    rr_2539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1207_inst_req_0); -- 
    rr_2553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1217_inst_req_0); -- 
    rr_2567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1227_inst_req_0); -- 
    rr_2581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1237_inst_req_0); -- 
    rr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => type_cast_1247_inst_req_0); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Sample/ra
      -- 
    ra_2498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_0, ack => convTranspose_CP_34_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	386 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	354 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Update/ca
      -- 
    ca_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_1, ack => convTranspose_CP_34_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	317 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Sample/ra
      -- 
    ra_2512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1187_inst_ack_0, ack => convTranspose_CP_34_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	386 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	351 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Update/ca
      -- 
    ca_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1187_inst_ack_1, ack => convTranspose_CP_34_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	317 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_sample_completed_
      -- CP-element group 322: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Sample/ra
      -- 
    ra_2526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_0, ack => convTranspose_CP_34_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	386 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	348 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_update_completed_
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Update/$exit
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Update/ca
      -- 
    ca_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_1, ack => convTranspose_CP_34_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	317 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Sample/ra
      -- 
    ra_2540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_0, ack => convTranspose_CP_34_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	386 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	345 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Update/ca
      -- 
    ca_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_1, ack => convTranspose_CP_34_elements(325)); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	317 
    -- CP-element group 326: successors 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_sample_completed_
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Sample/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Sample/ra
      -- 
    ra_2554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1217_inst_ack_0, ack => convTranspose_CP_34_elements(326)); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	386 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	342 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_update_completed_
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Update/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Update/ca
      -- 
    ca_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1217_inst_ack_1, ack => convTranspose_CP_34_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	317 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_sample_completed_
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Sample/ra
      -- 
    ra_2568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_0, ack => convTranspose_CP_34_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	386 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	339 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_update_completed_
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Update/ca
      -- 
    ca_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_1, ack => convTranspose_CP_34_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	317 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_sample_completed_
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Sample/ra
      -- 
    ra_2582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1237_inst_ack_0, ack => convTranspose_CP_34_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	386 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	336 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_update_completed_
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Update/ca
      -- 
    ca_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1237_inst_ack_1, ack => convTranspose_CP_34_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	317 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Sample/ra
      -- 
    ra_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_0, ack => convTranspose_CP_34_elements(332)); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	386 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Update/ca
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Sample/req
      -- 
    ca_2601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_1, ack => convTranspose_CP_34_elements(333)); -- 
    req_2609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(333), ack => WPIPE_ConvTranspose_output_pipe_1249_inst_req_0); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_sample_completed_
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_update_start_
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Sample/ack
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Update/req
      -- 
    ack_2610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1249_inst_ack_0, ack => convTranspose_CP_34_elements(334)); -- 
    req_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(334), ack => WPIPE_ConvTranspose_output_pipe_1249_inst_req_1); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1249_Update/ack
      -- 
    ack_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1249_inst_ack_1, ack => convTranspose_CP_34_elements(335)); -- 
    -- CP-element group 336:  join  transition  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	331 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Sample/req
      -- 
    req_2623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(336), ack => WPIPE_ConvTranspose_output_pipe_1252_inst_req_0); -- 
    convTranspose_cp_element_group_336: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_336"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(331) & convTranspose_CP_34_elements(335);
      gj_convTranspose_cp_element_group_336 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(336), clk => clk, reset => reset); --
    end block;
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_update_start_
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Update/req
      -- 
    ack_2624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1252_inst_ack_0, ack => convTranspose_CP_34_elements(337)); -- 
    req_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(337), ack => WPIPE_ConvTranspose_output_pipe_1252_inst_req_1); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1252_Update/ack
      -- 
    ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1252_inst_ack_1, ack => convTranspose_CP_34_elements(338)); -- 
    -- CP-element group 339:  join  transition  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	329 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Sample/req
      -- 
    req_2637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(339), ack => WPIPE_ConvTranspose_output_pipe_1255_inst_req_0); -- 
    convTranspose_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(329) & convTranspose_CP_34_elements(338);
      gj_convTranspose_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_update_start_
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Sample/ack
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Update/req
      -- 
    ack_2638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1255_inst_ack_0, ack => convTranspose_CP_34_elements(340)); -- 
    req_2642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(340), ack => WPIPE_ConvTranspose_output_pipe_1255_inst_req_1); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1255_Update/ack
      -- 
    ack_2643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1255_inst_ack_1, ack => convTranspose_CP_34_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	327 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Sample/req
      -- 
    req_2651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(342), ack => WPIPE_ConvTranspose_output_pipe_1258_inst_req_0); -- 
    convTranspose_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(327) & convTranspose_CP_34_elements(341);
      gj_convTranspose_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_update_start_
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Update/req
      -- 
    ack_2652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1258_inst_ack_0, ack => convTranspose_CP_34_elements(343)); -- 
    req_2656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(343), ack => WPIPE_ConvTranspose_output_pipe_1258_inst_req_1); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1258_Update/ack
      -- 
    ack_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1258_inst_ack_1, ack => convTranspose_CP_34_elements(344)); -- 
    -- CP-element group 345:  join  transition  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	325 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Sample/req
      -- 
    req_2665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(345), ack => WPIPE_ConvTranspose_output_pipe_1261_inst_req_0); -- 
    convTranspose_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(325) & convTranspose_CP_34_elements(344);
      gj_convTranspose_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_sample_completed_
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_update_start_
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Sample/ack
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Update/req
      -- 
    ack_2666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1261_inst_ack_0, ack => convTranspose_CP_34_elements(346)); -- 
    req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(346), ack => WPIPE_ConvTranspose_output_pipe_1261_inst_req_1); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_update_completed_
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1261_Update/ack
      -- 
    ack_2671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1261_inst_ack_1, ack => convTranspose_CP_34_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	323 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Sample/req
      -- 
    req_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(348), ack => WPIPE_ConvTranspose_output_pipe_1264_inst_req_0); -- 
    convTranspose_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(323) & convTranspose_CP_34_elements(347);
      gj_convTranspose_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  transition  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (6) 
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_update_start_
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Sample/ack
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Update/req
      -- 
    ack_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1264_inst_ack_0, ack => convTranspose_CP_34_elements(349)); -- 
    req_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(349), ack => WPIPE_ConvTranspose_output_pipe_1264_inst_req_1); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1264_Update/ack
      -- 
    ack_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1264_inst_ack_1, ack => convTranspose_CP_34_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	321 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Sample/req
      -- 
    req_2693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(351), ack => WPIPE_ConvTranspose_output_pipe_1267_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(321) & convTranspose_CP_34_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_update_start_
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Update/req
      -- 
    ack_2694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1267_inst_ack_0, ack => convTranspose_CP_34_elements(352)); -- 
    req_2698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(352), ack => WPIPE_ConvTranspose_output_pipe_1267_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1267_Update/ack
      -- 
    ack_2699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1267_inst_ack_1, ack => convTranspose_CP_34_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	319 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Sample/req
      -- 
    req_2707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(354), ack => WPIPE_ConvTranspose_output_pipe_1270_inst_req_0); -- 
    convTranspose_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(319) & convTranspose_CP_34_elements(353);
      gj_convTranspose_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (6) 
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_update_start_
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Sample/ack
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Update/req
      -- 
    ack_2708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1270_inst_ack_0, ack => convTranspose_CP_34_elements(355)); -- 
    req_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(355), ack => WPIPE_ConvTranspose_output_pipe_1270_inst_req_1); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/WPIPE_ConvTranspose_output_pipe_1270_Update/ack
      -- 
    ack_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1270_inst_ack_1, ack => convTranspose_CP_34_elements(356)); -- 
    -- CP-element group 357:  branch  join  transition  place  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	312 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (10) 
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283__exit__
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284__entry__
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/$exit
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284_dead_link/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284_eval_test/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284_eval_test/$exit
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284_eval_test/branch_req
      -- CP-element group 357: 	 branch_block_stmt_32/R_exitcond1_1285_place
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284_if_link/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/if_stmt_1284_else_link/$entry
      -- 
    branch_req_2721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(357), ack => if_stmt_1284_branch_req_0); -- 
    convTranspose_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(312) & convTranspose_CP_34_elements(356);
      gj_convTranspose_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  merge  transition  place  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	387 
    -- CP-element group 358:  members (13) 
      -- CP-element group 358: 	 branch_block_stmt_32/merge_stmt_1290__exit__
      -- CP-element group 358: 	 branch_block_stmt_32/forx_xend443x_xloopexit_forx_xend443
      -- CP-element group 358: 	 branch_block_stmt_32/forx_xend443x_xloopexit_forx_xend443_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/forx_xend443x_xloopexit_forx_xend443_PhiReq/$entry
      -- CP-element group 358: 	 branch_block_stmt_32/merge_stmt_1290_PhiReqMerge
      -- CP-element group 358: 	 branch_block_stmt_32/merge_stmt_1290_PhiAck/dummy
      -- CP-element group 358: 	 branch_block_stmt_32/merge_stmt_1290_PhiAck/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/merge_stmt_1290_PhiAck/$entry
      -- CP-element group 358: 	 branch_block_stmt_32/if_stmt_1284_if_link/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/if_stmt_1284_if_link/if_choice_transition
      -- CP-element group 358: 	 branch_block_stmt_32/forx_xbody370_forx_xend443x_xloopexit
      -- CP-element group 358: 	 branch_block_stmt_32/forx_xbody370_forx_xend443x_xloopexit_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/forx_xbody370_forx_xend443x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1284_branch_ack_1, ack => convTranspose_CP_34_elements(358)); -- 
    -- CP-element group 359:  fork  transition  place  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	382 
    -- CP-element group 359: 	383 
    -- CP-element group 359:  members (12) 
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Sample/rr
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Update/cr
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/if_stmt_1284_else_link/$exit
      -- CP-element group 359: 	 branch_block_stmt_32/if_stmt_1284_else_link/else_choice_transition
      -- CP-element group 359: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370
      -- 
    else_choice_transition_2730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1284_branch_ack_0, ack => convTranspose_CP_34_elements(359)); -- 
    rr_3005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(359), ack => type_cast_1162_inst_req_0); -- 
    cr_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(359), ack => type_cast_1162_inst_req_1); -- 
    -- CP-element group 360:  merge  branch  transition  place  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	120 
    -- CP-element group 360: 	165 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	121 
    -- CP-element group 360: 	122 
    -- CP-element group 360:  members (17) 
      -- CP-element group 360: 	 branch_block_stmt_32/merge_stmt_400__exit__
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_406__entry__
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_406__exit__
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407__entry__
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_406/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_406/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407_dead_link/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407_eval_test/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407_eval_test/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407_eval_test/branch_req
      -- CP-element group 360: 	 branch_block_stmt_32/R_cmp194452_408_place
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407_if_link/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/if_stmt_407_else_link/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/merge_stmt_400_PhiReqMerge
      -- CP-element group 360: 	 branch_block_stmt_32/merge_stmt_400_PhiAck/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/merge_stmt_400_PhiAck/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/merge_stmt_400_PhiAck/dummy
      -- 
    branch_req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(360), ack => if_stmt_407_branch_req_0); -- 
    convTranspose_CP_34_elements(360) <= OrReduce(convTranspose_CP_34_elements(120) & convTranspose_CP_34_elements(165));
    -- CP-element group 361:  transition  output  delay-element  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	124 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	365 
    -- CP-element group 361:  members (5) 
      -- CP-element group 361: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_451/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_455_konst_delay_trans
      -- CP-element group 361: 	 branch_block_stmt_32/bbx_xnph458_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_req
      -- 
    phi_stmt_451_req_2778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_451_req_2778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(361), ack => phi_stmt_451_req_0); -- 
    -- Element group convTranspose_CP_34_elements(361) is a control-delay.
    cp_element_361_delay: control_delay_element  generic map(name => " 361_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(124), ack => convTranspose_CP_34_elements(361), clk => clk, reset =>reset);
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	166 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Sample/ra
      -- 
    ra_2798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_0, ack => convTranspose_CP_34_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	166 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/Update/ca
      -- 
    ca_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_1, ack => convTranspose_CP_34_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (6) 
      -- CP-element group 364: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_sources/type_cast_457/SplitProtocol/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_451/phi_stmt_451_req
      -- 
    phi_stmt_451_req_2804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_451_req_2804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(364), ack => phi_stmt_451_req_1); -- 
    convTranspose_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(362) & convTranspose_CP_34_elements(363);
      gj_convTranspose_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  merge  transition  place  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	361 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (2) 
      -- CP-element group 365: 	 branch_block_stmt_32/merge_stmt_450_PhiReqMerge
      -- CP-element group 365: 	 branch_block_stmt_32/merge_stmt_450_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(365) <= OrReduce(convTranspose_CP_34_elements(361) & convTranspose_CP_34_elements(364));
    -- CP-element group 366:  fork  transition  place  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	125 
    -- CP-element group 366: 	126 
    -- CP-element group 366: 	128 
    -- CP-element group 366: 	129 
    -- CP-element group 366: 	132 
    -- CP-element group 366: 	136 
    -- CP-element group 366: 	140 
    -- CP-element group 366: 	144 
    -- CP-element group 366: 	148 
    -- CP-element group 366: 	152 
    -- CP-element group 366: 	156 
    -- CP-element group 366: 	160 
    -- CP-element group 366: 	163 
    -- CP-element group 366:  members (56) 
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_scale_1/scale_rename_ack
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/word_access_complete/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_scale_1/scale_rename_req
      -- CP-element group 366: 	 branch_block_stmt_32/merge_stmt_450__exit__
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613__entry__
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_scale_1/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_scale_1/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_resize_1/index_resize_ack
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_resize_1/index_resize_req
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_resize_1/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_resize_1/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_computed_1
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_scaled_1
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_index_resized_1
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_471_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Sample/rr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_556_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/RPIPE_ConvTranspose_input_pipe_467_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_574_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_502_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_520_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_complete/req
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/word_access_complete/word_0/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/addr_of_464_complete/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_592_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/ptr_deref_600_Update/word_access_complete/word_0/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Update/req
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_538_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Update/cr
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Sample/req
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/array_obj_ref_463_final_index_sum_regn_update_start
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_465_to_assign_stmt_613/type_cast_484_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/merge_stmt_450_PhiAck/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/merge_stmt_450_PhiAck/phi_stmt_451_ack
      -- 
    phi_stmt_451_ack_2809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_451_ack_0, ack => convTranspose_CP_34_elements(366)); -- 
    cr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_471_inst_req_1); -- 
    cr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_502_inst_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_556_inst_req_1); -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_574_inst_req_1); -- 
    cr_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_538_inst_req_1); -- 
    rr_1009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => RPIPE_ConvTranspose_input_pipe_467_inst_req_0); -- 
    cr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_520_inst_req_1); -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => addr_of_464_final_reg_req_1); -- 
    cr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_592_inst_req_1); -- 
    cr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => ptr_deref_600_store_0_req_1); -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => array_obj_ref_463_index_offset_req_1); -- 
    cr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => type_cast_484_inst_req_1); -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => array_obj_ref_463_index_offset_req_0); -- 
    -- CP-element group 367:  transition  output  delay-element  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	168 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	371 
    -- CP-element group 367:  members (5) 
      -- CP-element group 367: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_658/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_662_konst_delay_trans
      -- CP-element group 367: 	 branch_block_stmt_32/bbx_xnph454_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_req
      -- 
    phi_stmt_658_req_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_658_req_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(367), ack => phi_stmt_658_req_0); -- 
    -- Element group convTranspose_CP_34_elements(367) is a control-delay.
    cp_element_367_delay: control_delay_element  generic map(name => " 367_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(168), ack => convTranspose_CP_34_elements(367), clk => clk, reset =>reset);
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	210 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (2) 
      -- CP-element group 368: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Sample/ra
      -- 
    ra_2852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_0, ack => convTranspose_CP_34_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	210 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/Update/ca
      -- 
    ca_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_1, ack => convTranspose_CP_34_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_sources/type_cast_664/SplitProtocol/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_658/phi_stmt_658_req
      -- 
    phi_stmt_658_req_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_658_req_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(370), ack => phi_stmt_658_req_1); -- 
    convTranspose_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(368) & convTranspose_CP_34_elements(369);
      gj_convTranspose_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  merge  transition  place  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	367 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_32/merge_stmt_657_PhiReqMerge
      -- CP-element group 371: 	 branch_block_stmt_32/merge_stmt_657_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(371) <= OrReduce(convTranspose_CP_34_elements(367) & convTranspose_CP_34_elements(370));
    -- CP-element group 372:  fork  transition  place  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	207 
    -- CP-element group 372: 	204 
    -- CP-element group 372: 	169 
    -- CP-element group 372: 	170 
    -- CP-element group 372: 	172 
    -- CP-element group 372: 	173 
    -- CP-element group 372: 	176 
    -- CP-element group 372: 	180 
    -- CP-element group 372: 	184 
    -- CP-element group 372: 	188 
    -- CP-element group 372: 	192 
    -- CP-element group 372: 	196 
    -- CP-element group 372: 	200 
    -- CP-element group 372:  members (56) 
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_complete/req
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_691_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/merge_stmt_657__exit__
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820__entry__
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_resize_1/index_resize_ack
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_complete/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_resize_1/index_resize_req
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_resize_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_resize_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_computed_1
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_scaled_1
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_resized_1
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Sample/req
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/addr_of_671_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_update_start
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_scale_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Sample/rr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_scale_1/scale_rename_ack
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_678_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_scale_1/scale_rename_req
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_index_scale_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/array_obj_ref_670_final_index_sum_regn_Update/req
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/RPIPE_ConvTranspose_input_pipe_674_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_709_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_727_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_745_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_763_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_781_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/type_cast_799_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/word_access_complete/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/word_access_complete/word_0/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_672_to_assign_stmt_820/ptr_deref_807_Update/word_access_complete/word_0/cr
      -- CP-element group 372: 	 branch_block_stmt_32/merge_stmt_657_PhiAck/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/merge_stmt_657_PhiAck/phi_stmt_658_ack
      -- 
    phi_stmt_658_ack_2863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_658_ack_0, ack => convTranspose_CP_34_elements(372)); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_691_inst_req_1); -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => addr_of_671_final_reg_req_1); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => array_obj_ref_670_index_offset_req_0); -- 
    rr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => RPIPE_ConvTranspose_input_pipe_674_inst_req_0); -- 
    cr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_678_inst_req_1); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => array_obj_ref_670_index_offset_req_1); -- 
    cr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_709_inst_req_1); -- 
    cr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_727_inst_req_1); -- 
    cr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_745_inst_req_1); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_763_inst_req_1); -- 
    cr_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_781_inst_req_1); -- 
    cr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => type_cast_799_inst_req_1); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => ptr_deref_807_store_0_req_1); -- 
    -- CP-element group 373:  merge  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	209 
    -- CP-element group 373: 	122 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	211 
    -- CP-element group 373: 	212 
    -- CP-element group 373: 	213 
    -- CP-element group 373: 	214 
    -- CP-element group 373: 	215 
    -- CP-element group 373: 	216 
    -- CP-element group 373:  members (25) 
      -- CP-element group 373: 	 branch_block_stmt_32/merge_stmt_829__exit__
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857__entry__
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Sample/rr
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_832_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Sample/rr
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_836_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Sample/rr
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_833_to_assign_stmt_857/type_cast_840_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/merge_stmt_829_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_32/merge_stmt_829_PhiAck/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/merge_stmt_829_PhiAck/$exit
      -- CP-element group 373: 	 branch_block_stmt_32/merge_stmt_829_PhiAck/dummy
      -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_832_inst_req_0); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_832_inst_req_1); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_836_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_836_inst_req_1); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_840_inst_req_0); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_840_inst_req_1); -- 
    convTranspose_CP_34_elements(373) <= OrReduce(convTranspose_CP_34_elements(209) & convTranspose_CP_34_elements(122));
    -- CP-element group 374:  transition  output  delay-element  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	221 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	378 
    -- CP-element group 374:  members (5) 
      -- CP-element group 374: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_req
      -- CP-element group 374: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_906_konst_delay_trans
      -- CP-element group 374: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_902/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/bbx_xnph450_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/$exit
      -- 
    phi_stmt_902_req_2909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_902_req_2909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => phi_stmt_902_req_0); -- 
    -- Element group convTranspose_CP_34_elements(374) is a control-delay.
    cp_element_374_delay: control_delay_element  generic map(name => " 374_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(221), ack => convTranspose_CP_34_elements(374), clk => clk, reset =>reset);
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	230 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (2) 
      -- CP-element group 375: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Sample/ra
      -- CP-element group 375: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Sample/$exit
      -- 
    ra_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_0, ack => convTranspose_CP_34_elements(375)); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	230 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (2) 
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/Update/ca
      -- 
    ca_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_1, ack => convTranspose_CP_34_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/SplitProtocol/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_req
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_908/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_902/phi_stmt_902_sources/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- 
    phi_stmt_902_req_2935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_902_req_2935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => phi_stmt_902_req_1); -- 
    convTranspose_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(375) & convTranspose_CP_34_elements(376);
      gj_convTranspose_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  merge  transition  place  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	374 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_901_PhiAck/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_901_PhiReqMerge
      -- 
    convTranspose_CP_34_elements(378) <= OrReduce(convTranspose_CP_34_elements(374) & convTranspose_CP_34_elements(377));
    -- CP-element group 379:  fork  transition  place  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	227 
    -- CP-element group 379: 	222 
    -- CP-element group 379: 	223 
    -- CP-element group 379: 	225 
    -- CP-element group 379:  members (29) 
      -- CP-element group 379: 	 branch_block_stmt_32/merge_stmt_901__exit__
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932__entry__
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_update_start_
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_resized_1
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_scaled_1
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_computed_1
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_resize_1/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_resize_1/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_resize_1/index_resize_req
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_resize_1/index_resize_ack
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_scale_1/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_scale_1/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_scale_1/scale_rename_req
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_index_scale_1/scale_rename_ack
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_update_start
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Sample/req
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/array_obj_ref_914_final_index_sum_regn_Update/req
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_complete/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/addr_of_915_complete/req
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_update_start_
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/word_access_complete/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/word_access_complete/word_0/$entry
      -- CP-element group 379: 	 branch_block_stmt_32/assign_stmt_916_to_assign_stmt_932/ptr_deref_918_Update/word_access_complete/word_0/cr
      -- CP-element group 379: 	 branch_block_stmt_32/merge_stmt_901_PhiAck/phi_stmt_902_ack
      -- CP-element group 379: 	 branch_block_stmt_32/merge_stmt_901_PhiAck/$exit
      -- 
    phi_stmt_902_ack_2940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_902_ack_0, ack => convTranspose_CP_34_elements(379)); -- 
    req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(379), ack => array_obj_ref_914_index_offset_req_0); -- 
    req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(379), ack => array_obj_ref_914_index_offset_req_1); -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(379), ack => addr_of_915_final_reg_req_1); -- 
    cr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(379), ack => ptr_deref_918_store_0_req_1); -- 
    -- CP-element group 380:  merge  fork  transition  place  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	219 
    -- CP-element group 380: 	229 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	231 
    -- CP-element group 380: 	232 
    -- CP-element group 380: 	234 
    -- CP-element group 380:  members (16) 
      -- CP-element group 380: 	 branch_block_stmt_32/merge_stmt_941__exit__
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950__entry__
      -- CP-element group 380: 	 branch_block_stmt_32/merge_stmt_941_PhiReqMerge
      -- CP-element group 380: 	 branch_block_stmt_32/merge_stmt_941_PhiAck/$entry
      -- CP-element group 380: 	 branch_block_stmt_32/merge_stmt_941_PhiAck/$exit
      -- CP-element group 380: 	 branch_block_stmt_32/merge_stmt_941_PhiAck/dummy
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/$entry
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_update_start_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Sample/crr
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/call_stmt_944_Update/ccr
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_update_start_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_944_to_assign_stmt_950/type_cast_949_Update/cr
      -- 
    crr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(380), ack => call_stmt_944_call_req_0); -- 
    ccr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(380), ack => call_stmt_944_call_req_1); -- 
    cr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(380), ack => type_cast_949_inst_req_1); -- 
    convTranspose_CP_34_elements(380) <= OrReduce(convTranspose_CP_34_elements(219) & convTranspose_CP_34_elements(229));
    -- CP-element group 381:  transition  output  delay-element  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	311 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	385 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_req
      -- CP-element group 381: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1160_konst_delay_trans
      -- CP-element group 381: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/phi_stmt_1156/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/bbx_xnph_forx_xbody370_PhiReq/$exit
      -- 
    phi_stmt_1156_req_2986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1156_req_2986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(381), ack => phi_stmt_1156_req_0); -- 
    -- Element group convTranspose_CP_34_elements(381) is a control-delay.
    cp_element_381_delay: control_delay_element  generic map(name => " 381_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(311), ack => convTranspose_CP_34_elements(381), clk => clk, reset =>reset);
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	359 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (2) 
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Sample/ra
      -- 
    ra_3006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_0, ack => convTranspose_CP_34_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	359 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (2) 
      -- CP-element group 383: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/Update/ca
      -- 
    ca_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_1, ack => convTranspose_CP_34_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/SplitProtocol/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/type_cast_1162/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_sources/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/phi_stmt_1156_req
      -- CP-element group 384: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/phi_stmt_1156/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/forx_xbody370_forx_xbody370_PhiReq/$exit
      -- 
    phi_stmt_1156_req_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1156_req_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(384), ack => phi_stmt_1156_req_1); -- 
    convTranspose_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(382) & convTranspose_CP_34_elements(383);
      gj_convTranspose_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  merge  transition  place  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	381 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (2) 
      -- CP-element group 385: 	 branch_block_stmt_32/merge_stmt_1155_PhiReqMerge
      -- CP-element group 385: 	 branch_block_stmt_32/merge_stmt_1155_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(385) <= OrReduce(convTranspose_CP_34_elements(381) & convTranspose_CP_34_elements(384));
    -- CP-element group 386:  fork  transition  place  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	312 
    -- CP-element group 386: 	313 
    -- CP-element group 386: 	315 
    -- CP-element group 386: 	317 
    -- CP-element group 386: 	319 
    -- CP-element group 386: 	321 
    -- CP-element group 386: 	323 
    -- CP-element group 386: 	325 
    -- CP-element group 386: 	327 
    -- CP-element group 386: 	329 
    -- CP-element group 386: 	331 
    -- CP-element group 386: 	333 
    -- CP-element group 386:  members (53) 
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_scale_1/$exit
      -- CP-element group 386: 	 branch_block_stmt_32/merge_stmt_1155__exit__
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283__entry__
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Sample/req
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_scale_1/scale_rename_req
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_scale_1/scale_rename_ack
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_resize_1/index_resize_req
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_scale_1/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Update/req
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_resize_1/$exit
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_update_start
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_resize_1/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_final_index_sum_regn_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_computed_1
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_resize_1/index_resize_ack
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_scaled_1
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/array_obj_ref_1168_index_resized_1
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_complete/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/addr_of_1169_complete/req
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/word_access_complete/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/word_access_complete/word_0/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/ptr_deref_1173_Update/word_access_complete/word_0/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1177_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1187_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1197_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1207_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1217_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1227_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1237_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/assign_stmt_1170_to_assign_stmt_1283/type_cast_1247_Update/cr
      -- CP-element group 386: 	 branch_block_stmt_32/merge_stmt_1155_PhiAck/phi_stmt_1156_ack
      -- CP-element group 386: 	 branch_block_stmt_32/merge_stmt_1155_PhiAck/$exit
      -- 
    phi_stmt_1156_ack_3017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1156_ack_0, ack => convTranspose_CP_34_elements(386)); -- 
    req_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => array_obj_ref_1168_index_offset_req_0); -- 
    req_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => array_obj_ref_1168_index_offset_req_1); -- 
    req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => addr_of_1169_final_reg_req_1); -- 
    cr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => ptr_deref_1173_load_0_req_1); -- 
    cr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1177_inst_req_1); -- 
    cr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1187_inst_req_1); -- 
    cr_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1197_inst_req_1); -- 
    cr_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1207_inst_req_1); -- 
    cr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1217_inst_req_1); -- 
    cr_2572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1227_inst_req_1); -- 
    cr_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1237_inst_req_1); -- 
    cr_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(386), ack => type_cast_1247_inst_req_1); -- 
    -- CP-element group 387:  merge  transition  place  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	309 
    -- CP-element group 387: 	358 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (16) 
      -- CP-element group 387: 	 $exit
      -- CP-element group 387: 	 branch_block_stmt_32/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1292__exit__
      -- CP-element group 387: 	 branch_block_stmt_32/return__
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1294__exit__
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1292_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1292_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1294_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1294_PhiAck/dummy
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1294_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1292_PhiReqMerge
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1292_PhiAck/dummy
      -- CP-element group 387: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 387: 	 branch_block_stmt_32/merge_stmt_1294_PhiReqMerge
      -- CP-element group 387: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- 
    convTranspose_CP_34_elements(387) <= OrReduce(convTranspose_CP_34_elements(309) & convTranspose_CP_34_elements(358));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar468_913_resized : std_logic_vector(13 downto 0);
    signal R_indvar468_913_scaled : std_logic_vector(13 downto 0);
    signal R_indvar482_669_resized : std_logic_vector(10 downto 0);
    signal R_indvar482_669_scaled : std_logic_vector(10 downto 0);
    signal R_indvar498_462_resized : std_logic_vector(13 downto 0);
    signal R_indvar498_462_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1167_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1167_scaled : std_logic_vector(13 downto 0);
    signal add108_310 : std_logic_vector(15 downto 0);
    signal add117_335 : std_logic_vector(15 downto 0);
    signal add126_360 : std_logic_vector(15 downto 0);
    signal add12_82 : std_logic_vector(15 downto 0);
    signal add135_385 : std_logic_vector(15 downto 0);
    signal add150_490 : std_logic_vector(63 downto 0);
    signal add156_508 : std_logic_vector(63 downto 0);
    signal add162_526 : std_logic_vector(63 downto 0);
    signal add168_544 : std_logic_vector(63 downto 0);
    signal add174_562 : std_logic_vector(63 downto 0);
    signal add180_580 : std_logic_vector(63 downto 0);
    signal add186_598 : std_logic_vector(63 downto 0);
    signal add206_697 : std_logic_vector(63 downto 0);
    signal add212_715 : std_logic_vector(63 downto 0);
    signal add218_733 : std_logic_vector(63 downto 0);
    signal add21_107 : std_logic_vector(15 downto 0);
    signal add224_751 : std_logic_vector(63 downto 0);
    signal add230_769 : std_logic_vector(63 downto 0);
    signal add236_787 : std_logic_vector(63 downto 0);
    signal add242_805 : std_logic_vector(63 downto 0);
    signal add30_132 : std_logic_vector(15 downto 0);
    signal add39_157 : std_logic_vector(15 downto 0);
    signal add48_182 : std_logic_vector(15 downto 0);
    signal add57_207 : std_logic_vector(15 downto 0);
    signal add99_285 : std_logic_vector(15 downto 0);
    signal add_57 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1168_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1168_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1168_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1168_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1168_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1168_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_463_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_463_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_463_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_463_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_463_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_463_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_670_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_670_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_670_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_670_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_670_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_670_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_914_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_914_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_914_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_914_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_914_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_914_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_672 : std_logic_vector(31 downto 0);
    signal arrayidx269_916 : std_logic_vector(31 downto 0);
    signal arrayidx375_1170 : std_logic_vector(31 downto 0);
    signal arrayidx_465 : std_logic_vector(31 downto 0);
    signal call101_288 : std_logic_vector(7 downto 0);
    signal call106_301 : std_logic_vector(7 downto 0);
    signal call10_73 : std_logic_vector(7 downto 0);
    signal call110_313 : std_logic_vector(7 downto 0);
    signal call115_326 : std_logic_vector(7 downto 0);
    signal call119_338 : std_logic_vector(7 downto 0);
    signal call124_351 : std_logic_vector(7 downto 0);
    signal call128_363 : std_logic_vector(7 downto 0);
    signal call133_376 : std_logic_vector(7 downto 0);
    signal call143_468 : std_logic_vector(7 downto 0);
    signal call147_481 : std_logic_vector(7 downto 0);
    signal call14_85 : std_logic_vector(7 downto 0);
    signal call153_499 : std_logic_vector(7 downto 0);
    signal call159_517 : std_logic_vector(7 downto 0);
    signal call165_535 : std_logic_vector(7 downto 0);
    signal call171_553 : std_logic_vector(7 downto 0);
    signal call177_571 : std_logic_vector(7 downto 0);
    signal call183_589 : std_logic_vector(7 downto 0);
    signal call199_675 : std_logic_vector(7 downto 0);
    signal call19_98 : std_logic_vector(7 downto 0);
    signal call203_688 : std_logic_vector(7 downto 0);
    signal call209_706 : std_logic_vector(7 downto 0);
    signal call215_724 : std_logic_vector(7 downto 0);
    signal call221_742 : std_logic_vector(7 downto 0);
    signal call227_760 : std_logic_vector(7 downto 0);
    signal call233_778 : std_logic_vector(7 downto 0);
    signal call239_796 : std_logic_vector(7 downto 0);
    signal call23_110 : std_logic_vector(7 downto 0);
    signal call275_944 : std_logic_vector(63 downto 0);
    signal call28_123 : std_logic_vector(7 downto 0);
    signal call295_999 : std_logic_vector(15 downto 0);
    signal call297_1002 : std_logic_vector(63 downto 0);
    signal call2_48 : std_logic_vector(7 downto 0);
    signal call32_135 : std_logic_vector(7 downto 0);
    signal call37_148 : std_logic_vector(7 downto 0);
    signal call41_160 : std_logic_vector(7 downto 0);
    signal call46_173 : std_logic_vector(7 downto 0);
    signal call50_185 : std_logic_vector(7 downto 0);
    signal call55_198 : std_logic_vector(7 downto 0);
    signal call5_60 : std_logic_vector(7 downto 0);
    signal call92_263 : std_logic_vector(7 downto 0);
    signal call97_276 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp194452_406 : std_logic_vector(0 downto 0);
    signal cmp264448_857 : std_logic_vector(0 downto 0);
    signal cmp456_391 : std_logic_vector(0 downto 0);
    signal conv104_292 : std_logic_vector(15 downto 0);
    signal conv107_305 : std_logic_vector(15 downto 0);
    signal conv113_317 : std_logic_vector(15 downto 0);
    signal conv116_330 : std_logic_vector(15 downto 0);
    signal conv11_77 : std_logic_vector(15 downto 0);
    signal conv122_342 : std_logic_vector(15 downto 0);
    signal conv125_355 : std_logic_vector(15 downto 0);
    signal conv131_367 : std_logic_vector(15 downto 0);
    signal conv134_380 : std_logic_vector(15 downto 0);
    signal conv144_472 : std_logic_vector(63 downto 0);
    signal conv149_485 : std_logic_vector(63 downto 0);
    signal conv155_503 : std_logic_vector(63 downto 0);
    signal conv161_521 : std_logic_vector(63 downto 0);
    signal conv167_539 : std_logic_vector(63 downto 0);
    signal conv173_557 : std_logic_vector(63 downto 0);
    signal conv179_575 : std_logic_vector(63 downto 0);
    signal conv17_89 : std_logic_vector(15 downto 0);
    signal conv185_593 : std_logic_vector(63 downto 0);
    signal conv1_39 : std_logic_vector(15 downto 0);
    signal conv200_679 : std_logic_vector(63 downto 0);
    signal conv205_692 : std_logic_vector(63 downto 0);
    signal conv20_102 : std_logic_vector(15 downto 0);
    signal conv211_710 : std_logic_vector(63 downto 0);
    signal conv217_728 : std_logic_vector(63 downto 0);
    signal conv223_746 : std_logic_vector(63 downto 0);
    signal conv229_764 : std_logic_vector(63 downto 0);
    signal conv235_782 : std_logic_vector(63 downto 0);
    signal conv241_800 : std_logic_vector(63 downto 0);
    signal conv253_833 : std_logic_vector(31 downto 0);
    signal conv255_837 : std_logic_vector(31 downto 0);
    signal conv258_841 : std_logic_vector(31 downto 0);
    signal conv26_114 : std_logic_vector(15 downto 0);
    signal conv276_950 : std_logic_vector(63 downto 0);
    signal conv298_1007 : std_logic_vector(63 downto 0);
    signal conv29_127 : std_logic_vector(15 downto 0);
    signal conv304_1016 : std_logic_vector(7 downto 0);
    signal conv310_1026 : std_logic_vector(7 downto 0);
    signal conv316_1036 : std_logic_vector(7 downto 0);
    signal conv322_1046 : std_logic_vector(7 downto 0);
    signal conv328_1056 : std_logic_vector(7 downto 0);
    signal conv334_1066 : std_logic_vector(7 downto 0);
    signal conv340_1076 : std_logic_vector(7 downto 0);
    signal conv346_1086 : std_logic_vector(7 downto 0);
    signal conv35_139 : std_logic_vector(15 downto 0);
    signal conv380_1178 : std_logic_vector(7 downto 0);
    signal conv386_1188 : std_logic_vector(7 downto 0);
    signal conv38_152 : std_logic_vector(15 downto 0);
    signal conv392_1198 : std_logic_vector(7 downto 0);
    signal conv398_1208 : std_logic_vector(7 downto 0);
    signal conv3_52 : std_logic_vector(15 downto 0);
    signal conv404_1218 : std_logic_vector(7 downto 0);
    signal conv410_1228 : std_logic_vector(7 downto 0);
    signal conv416_1238 : std_logic_vector(7 downto 0);
    signal conv422_1248 : std_logic_vector(7 downto 0);
    signal conv44_164 : std_logic_vector(15 downto 0);
    signal conv47_177 : std_logic_vector(15 downto 0);
    signal conv53_189 : std_logic_vector(15 downto 0);
    signal conv56_202 : std_logic_vector(15 downto 0);
    signal conv61_211 : std_logic_vector(31 downto 0);
    signal conv63_215 : std_logic_vector(31 downto 0);
    signal conv65_219 : std_logic_vector(31 downto 0);
    signal conv82_233 : std_logic_vector(31 downto 0);
    signal conv84_237 : std_logic_vector(31 downto 0);
    signal conv87_241 : std_logic_vector(31 downto 0);
    signal conv8_64 : std_logic_vector(15 downto 0);
    signal conv90_245 : std_logic_vector(31 downto 0);
    signal conv95_267 : std_logic_vector(15 downto 0);
    signal conv98_280 : std_logic_vector(15 downto 0);
    signal exitcond1_1283 : std_logic_vector(0 downto 0);
    signal exitcond2_820 : std_logic_vector(0 downto 0);
    signal exitcond3_613 : std_logic_vector(0 downto 0);
    signal exitcond_932 : std_logic_vector(0 downto 0);
    signal iNsTr_108_1140 : std_logic_vector(63 downto 0);
    signal iNsTr_25_435 : std_logic_vector(63 downto 0);
    signal iNsTr_38_642 : std_logic_vector(63 downto 0);
    signal iNsTr_52_886 : std_logic_vector(63 downto 0);
    signal indvar468_902 : std_logic_vector(63 downto 0);
    signal indvar482_658 : std_logic_vector(63 downto 0);
    signal indvar498_451 : std_logic_vector(63 downto 0);
    signal indvar_1156 : std_logic_vector(63 downto 0);
    signal indvarx_xnext469_927 : std_logic_vector(63 downto 0);
    signal indvarx_xnext483_815 : std_logic_vector(63 downto 0);
    signal indvarx_xnext499_608 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1278 : std_logic_vector(63 downto 0);
    signal mul256_846 : std_logic_vector(31 downto 0);
    signal mul259_851 : std_logic_vector(31 downto 0);
    signal mul66_229 : std_logic_vector(31 downto 0);
    signal mul85_250 : std_logic_vector(31 downto 0);
    signal mul88_255 : std_logic_vector(31 downto 0);
    signal mul91_260 : std_logic_vector(31 downto 0);
    signal mul_224 : std_logic_vector(31 downto 0);
    signal ptr_deref_1173_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1173_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1173_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1173_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1173_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_600_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_600_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_600_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_600_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_600_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_600_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_807_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_807_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_807_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_807_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_807_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_807_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_918_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_918_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_918_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_918_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_918_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_918_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_298 : std_logic_vector(15 downto 0);
    signal shl114_323 : std_logic_vector(15 downto 0);
    signal shl123_348 : std_logic_vector(15 downto 0);
    signal shl132_373 : std_logic_vector(15 downto 0);
    signal shl146_478 : std_logic_vector(63 downto 0);
    signal shl152_496 : std_logic_vector(63 downto 0);
    signal shl158_514 : std_logic_vector(63 downto 0);
    signal shl164_532 : std_logic_vector(63 downto 0);
    signal shl170_550 : std_logic_vector(63 downto 0);
    signal shl176_568 : std_logic_vector(63 downto 0);
    signal shl182_586 : std_logic_vector(63 downto 0);
    signal shl18_95 : std_logic_vector(15 downto 0);
    signal shl202_685 : std_logic_vector(63 downto 0);
    signal shl208_703 : std_logic_vector(63 downto 0);
    signal shl214_721 : std_logic_vector(63 downto 0);
    signal shl220_739 : std_logic_vector(63 downto 0);
    signal shl226_757 : std_logic_vector(63 downto 0);
    signal shl232_775 : std_logic_vector(63 downto 0);
    signal shl238_793 : std_logic_vector(63 downto 0);
    signal shl27_120 : std_logic_vector(15 downto 0);
    signal shl36_145 : std_logic_vector(15 downto 0);
    signal shl45_170 : std_logic_vector(15 downto 0);
    signal shl54_195 : std_logic_vector(15 downto 0);
    signal shl96_273 : std_logic_vector(15 downto 0);
    signal shl9_70 : std_logic_vector(15 downto 0);
    signal shl_45 : std_logic_vector(15 downto 0);
    signal shr307_1022 : std_logic_vector(63 downto 0);
    signal shr313_1032 : std_logic_vector(63 downto 0);
    signal shr319_1042 : std_logic_vector(63 downto 0);
    signal shr325_1052 : std_logic_vector(63 downto 0);
    signal shr331_1062 : std_logic_vector(63 downto 0);
    signal shr337_1072 : std_logic_vector(63 downto 0);
    signal shr343_1082 : std_logic_vector(63 downto 0);
    signal shr383_1184 : std_logic_vector(63 downto 0);
    signal shr389_1194 : std_logic_vector(63 downto 0);
    signal shr395_1204 : std_logic_vector(63 downto 0);
    signal shr401_1214 : std_logic_vector(63 downto 0);
    signal shr407_1224 : std_logic_vector(63 downto 0);
    signal shr413_1234 : std_logic_vector(63 downto 0);
    signal shr419_1244 : std_logic_vector(63 downto 0);
    signal sub_1012 : std_logic_vector(63 downto 0);
    signal tmp376_1174 : std_logic_vector(63 downto 0);
    signal tmp463_1124 : std_logic_vector(31 downto 0);
    signal tmp463x_xop_1136 : std_logic_vector(31 downto 0);
    signal tmp464_1130 : std_logic_vector(0 downto 0);
    signal tmp467_1153 : std_logic_vector(63 downto 0);
    signal tmp475_870 : std_logic_vector(31 downto 0);
    signal tmp475x_xop_882 : std_logic_vector(31 downto 0);
    signal tmp476_876 : std_logic_vector(0 downto 0);
    signal tmp480_899 : std_logic_vector(63 downto 0);
    signal tmp491_626 : std_logic_vector(31 downto 0);
    signal tmp491x_xop_638 : std_logic_vector(31 downto 0);
    signal tmp492_632 : std_logic_vector(0 downto 0);
    signal tmp496_655 : std_logic_vector(63 downto 0);
    signal tmp505_419 : std_logic_vector(31 downto 0);
    signal tmp505x_xop_431 : std_logic_vector(31 downto 0);
    signal tmp506_425 : std_logic_vector(0 downto 0);
    signal tmp510_448 : std_logic_vector(63 downto 0);
    signal type_cast_1005_wire : std_logic_vector(63 downto 0);
    signal type_cast_1020_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1040_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1050_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1060_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1070_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1122_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1128_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1134_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1151_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1160_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1162_wire : std_logic_vector(63 downto 0);
    signal type_cast_1182_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1192_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1212_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1222_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1232_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1242_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_271_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_321_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_371_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_389_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_404_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_417_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_423_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_439_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_43_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_455_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_457_wire : std_logic_vector(63 downto 0);
    signal type_cast_476_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_630_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_646_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_653_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_662_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_664_wire : std_logic_vector(63 downto 0);
    signal type_cast_683_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_701_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_737_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_791_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_813_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_855_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_880_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_925_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_948_wire : std_logic_vector(63 downto 0);
    signal type_cast_981_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_985_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop512_892 : std_logic_vector(63 downto 0);
    signal xx_xop513_648 : std_logic_vector(63 downto 0);
    signal xx_xop514_441 : std_logic_vector(63 downto 0);
    signal xx_xop_1146 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1168_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1168_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1168_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1168_resized_base_address <= "00000000000000";
    array_obj_ref_463_constant_part_of_offset <= "00000000000000";
    array_obj_ref_463_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_463_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_463_resized_base_address <= "00000000000000";
    array_obj_ref_670_constant_part_of_offset <= "00000100010";
    array_obj_ref_670_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_670_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_670_resized_base_address <= "00000000000";
    array_obj_ref_914_constant_part_of_offset <= "00000000000000";
    array_obj_ref_914_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_914_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_914_resized_base_address <= "00000000000000";
    ptr_deref_1173_word_offset_0 <= "00000000000000";
    ptr_deref_600_word_offset_0 <= "00000000000000";
    ptr_deref_807_word_offset_0 <= "00000000000";
    ptr_deref_918_word_offset_0 <= "00000000000000";
    type_cast_1020_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1040_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1050_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1060_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1070_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1080_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1122_wire_constant <= "00000000000000000000000000000010";
    type_cast_1128_wire_constant <= "00000000000000000000000000000001";
    type_cast_1134_wire_constant <= "11111111111111111111111111111111";
    type_cast_1144_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1151_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1160_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1182_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_118_wire_constant <= "0000000000001000";
    type_cast_1192_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1202_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1212_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1232_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1242_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1276_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_143_wire_constant <= "0000000000001000";
    type_cast_168_wire_constant <= "0000000000001000";
    type_cast_193_wire_constant <= "0000000000001000";
    type_cast_271_wire_constant <= "0000000000001000";
    type_cast_296_wire_constant <= "0000000000001000";
    type_cast_321_wire_constant <= "0000000000001000";
    type_cast_346_wire_constant <= "0000000000001000";
    type_cast_371_wire_constant <= "0000000000001000";
    type_cast_389_wire_constant <= "00000000000000000000000000000011";
    type_cast_404_wire_constant <= "00000000000000000000000000000011";
    type_cast_417_wire_constant <= "00000000000000000000000000000010";
    type_cast_423_wire_constant <= "00000000000000000000000000000001";
    type_cast_429_wire_constant <= "11111111111111111111111111111111";
    type_cast_439_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_43_wire_constant <= "0000000000001000";
    type_cast_446_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_476_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_494_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_584_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_606_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_624_wire_constant <= "00000000000000000000000000000010";
    type_cast_630_wire_constant <= "00000000000000000000000000000001";
    type_cast_636_wire_constant <= "11111111111111111111111111111111";
    type_cast_646_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_653_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_662_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_683_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_68_wire_constant <= "0000000000001000";
    type_cast_701_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_737_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_791_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_813_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_855_wire_constant <= "00000000000000000000000000000011";
    type_cast_868_wire_constant <= "00000000000000000000000000000010";
    type_cast_874_wire_constant <= "00000000000000000000000000000001";
    type_cast_880_wire_constant <= "11111111111111111111111111111111";
    type_cast_890_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_897_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_906_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_925_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_93_wire_constant <= "0000000000001000";
    type_cast_981_wire_constant <= "0000000000000000";
    type_cast_985_wire_constant <= "0000000000000000";
    phi_stmt_1156: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1160_wire_constant & type_cast_1162_wire;
      req <= phi_stmt_1156_req_0 & phi_stmt_1156_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1156",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1156_ack_0,
          idata => idata,
          odata => indvar_1156,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1156
    phi_stmt_451: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_455_wire_constant & type_cast_457_wire;
      req <= phi_stmt_451_req_0 & phi_stmt_451_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_451",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_451_ack_0,
          idata => idata,
          odata => indvar498_451,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_451
    phi_stmt_658: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_662_wire_constant & type_cast_664_wire;
      req <= phi_stmt_658_req_0 & phi_stmt_658_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_658",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_658_ack_0,
          idata => idata,
          odata => indvar482_658,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_658
    phi_stmt_902: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_906_wire_constant & type_cast_908_wire;
      req <= phi_stmt_902_req_0 & phi_stmt_902_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_902",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_902_ack_0,
          idata => idata,
          odata => indvar468_902,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_902
    -- flow-through select operator MUX_1152_inst
    tmp467_1153 <= xx_xop_1146 when (tmp464_1130(0) /=  '0') else type_cast_1151_wire_constant;
    -- flow-through select operator MUX_447_inst
    tmp510_448 <= xx_xop514_441 when (tmp506_425(0) /=  '0') else type_cast_446_wire_constant;
    -- flow-through select operator MUX_654_inst
    tmp496_655 <= xx_xop513_648 when (tmp492_632(0) /=  '0') else type_cast_653_wire_constant;
    -- flow-through select operator MUX_898_inst
    tmp480_899 <= xx_xop512_892 when (tmp476_876(0) /=  '0') else type_cast_897_wire_constant;
    addr_of_1169_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1169_final_reg_req_0;
      addr_of_1169_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1169_final_reg_req_1;
      addr_of_1169_final_reg_ack_1<= rack(0);
      addr_of_1169_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1169_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1168_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx375_1170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_464_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_464_final_reg_req_0;
      addr_of_464_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_464_final_reg_req_1;
      addr_of_464_final_reg_ack_1<= rack(0);
      addr_of_464_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_464_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_463_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_465,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_671_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_671_final_reg_req_0;
      addr_of_671_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_671_final_reg_req_1;
      addr_of_671_final_reg_ack_1<= rack(0);
      addr_of_671_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_671_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_670_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_915_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_915_final_reg_req_0;
      addr_of_915_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_915_final_reg_req_1;
      addr_of_915_final_reg_ack_1<= rack(0);
      addr_of_915_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_915_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_914_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1006_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1006_inst_req_0;
      type_cast_1006_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1006_inst_req_1;
      type_cast_1006_inst_ack_1<= rack(0);
      type_cast_1006_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1006_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1005_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_1007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1015_inst_req_0;
      type_cast_1015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1015_inst_req_1;
      type_cast_1015_inst_ack_1<= rack(0);
      type_cast_1015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_1016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_101_inst_req_0;
      type_cast_101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_101_inst_req_1;
      type_cast_101_inst_ack_1<= rack(0);
      type_cast_101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1025_inst_req_0;
      type_cast_1025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1025_inst_req_1;
      type_cast_1025_inst_ack_1<= rack(0);
      type_cast_1025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr307_1022,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv310_1026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1035_inst_req_0;
      type_cast_1035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1035_inst_req_1;
      type_cast_1035_inst_ack_1<= rack(0);
      type_cast_1035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr313_1032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv316_1036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1045_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1045_inst_req_0;
      type_cast_1045_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1045_inst_req_1;
      type_cast_1045_inst_ack_1<= rack(0);
      type_cast_1045_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1045_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr319_1042,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1046,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr325_1052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv328_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1065_inst_req_0;
      type_cast_1065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1065_inst_req_1;
      type_cast_1065_inst_ack_1<= rack(0);
      type_cast_1065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr331_1062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv334_1066,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1075_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1075_inst_req_0;
      type_cast_1075_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1075_inst_req_1;
      type_cast_1075_inst_ack_1<= rack(0);
      type_cast_1075_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1075_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr337_1072,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv340_1076,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1085_inst_req_0;
      type_cast_1085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1085_inst_req_1;
      type_cast_1085_inst_ack_1<= rack(0);
      type_cast_1085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr343_1082,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv346_1086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1139_inst_req_0;
      type_cast_1139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1139_inst_req_1;
      type_cast_1139_inst_ack_1<= rack(0);
      type_cast_1139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp463x_xop_1136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_108_1140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1162_inst_req_0;
      type_cast_1162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1162_inst_req_1;
      type_cast_1162_inst_ack_1<= rack(0);
      type_cast_1162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1278,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1162_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1177_inst_req_0;
      type_cast_1177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1177_inst_req_1;
      type_cast_1177_inst_ack_1<= rack(0);
      type_cast_1177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp376_1174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv380_1178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1187_inst_req_0;
      type_cast_1187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1187_inst_req_1;
      type_cast_1187_inst_ack_1<= rack(0);
      type_cast_1187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr383_1184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv386_1188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1197_inst_req_0;
      type_cast_1197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1197_inst_req_1;
      type_cast_1197_inst_ack_1<= rack(0);
      type_cast_1197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr389_1194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv392_1198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1207_inst_req_0;
      type_cast_1207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1207_inst_req_1;
      type_cast_1207_inst_ack_1<= rack(0);
      type_cast_1207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr395_1204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv398_1208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1217_inst_req_0;
      type_cast_1217_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1217_inst_req_1;
      type_cast_1217_inst_ack_1<= rack(0);
      type_cast_1217_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1217_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr401_1214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv404_1218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1227_inst_req_0;
      type_cast_1227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1227_inst_req_1;
      type_cast_1227_inst_ack_1<= rack(0);
      type_cast_1227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr407_1224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv410_1228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1237_inst_req_0;
      type_cast_1237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1237_inst_req_1;
      type_cast_1237_inst_ack_1<= rack(0);
      type_cast_1237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr413_1234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv416_1238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1247_inst_req_0;
      type_cast_1247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1247_inst_req_1;
      type_cast_1247_inst_ack_1<= rack(0);
      type_cast_1247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr419_1244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv422_1248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_188_inst_req_0;
      type_cast_188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_188_inst_req_1;
      type_cast_188_inst_ack_1<= rack(0);
      type_cast_188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_210_inst_req_0;
      type_cast_210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_210_inst_req_1;
      type_cast_210_inst_ack_1<= rack(0);
      type_cast_210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_57,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_82,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_218_inst_req_0;
      type_cast_218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_218_inst_req_1;
      type_cast_218_inst_ack_1<= rack(0);
      type_cast_218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_232_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_232_inst_req_0;
      type_cast_232_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_232_inst_req_1;
      type_cast_232_inst_ack_1<= rack(0);
      type_cast_232_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_232_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_233,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_236_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_236_inst_req_0;
      type_cast_236_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_236_inst_req_1;
      type_cast_236_inst_ack_1<= rack(0);
      type_cast_236_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_236_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_237,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_240_inst_req_0;
      type_cast_240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_240_inst_req_1;
      type_cast_240_inst_ack_1<= rack(0);
      type_cast_240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_244_inst_req_0;
      type_cast_244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_244_inst_req_1;
      type_cast_244_inst_ack_1<= rack(0);
      type_cast_244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_245,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_266_inst_req_0;
      type_cast_266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_266_inst_req_1;
      type_cast_266_inst_ack_1<= rack(0);
      type_cast_266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_279_inst_req_0;
      type_cast_279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_279_inst_req_1;
      type_cast_279_inst_ack_1<= rack(0);
      type_cast_279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_291_inst_req_0;
      type_cast_291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_291_inst_req_1;
      type_cast_291_inst_ack_1<= rack(0);
      type_cast_291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_304_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_304_inst_req_0;
      type_cast_304_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_304_inst_req_1;
      type_cast_304_inst_ack_1<= rack(0);
      type_cast_304_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_304_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_316_inst_req_0;
      type_cast_316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_316_inst_req_1;
      type_cast_316_inst_ack_1<= rack(0);
      type_cast_316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_329_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_329_inst_req_0;
      type_cast_329_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_329_inst_req_1;
      type_cast_329_inst_ack_1<= rack(0);
      type_cast_329_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_329_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_326,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_330,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_341_inst_req_0;
      type_cast_341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_341_inst_req_1;
      type_cast_341_inst_ack_1<= rack(0);
      type_cast_341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_354_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_354_inst_req_0;
      type_cast_354_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_354_inst_req_1;
      type_cast_354_inst_ack_1<= rack(0);
      type_cast_354_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_354_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_351,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_355,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_366_inst_req_0;
      type_cast_366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_366_inst_req_1;
      type_cast_366_inst_ack_1<= rack(0);
      type_cast_366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_379_inst_req_0;
      type_cast_379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_379_inst_req_1;
      type_cast_379_inst_ack_1<= rack(0);
      type_cast_379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_379_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_380,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_434_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_434_inst_req_0;
      type_cast_434_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_434_inst_req_1;
      type_cast_434_inst_ack_1<= rack(0);
      type_cast_434_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_434_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp505x_xop_431,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_25_435,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_457_inst_req_0;
      type_cast_457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_457_inst_req_1;
      type_cast_457_inst_ack_1<= rack(0);
      type_cast_457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext499_608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_457_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_471_inst_req_0;
      type_cast_471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_471_inst_req_1;
      type_cast_471_inst_ack_1<= rack(0);
      type_cast_471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_468,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_484_inst_req_0;
      type_cast_484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_484_inst_req_1;
      type_cast_484_inst_ack_1<= rack(0);
      type_cast_484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_481,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_502_inst_req_0;
      type_cast_502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_502_inst_req_1;
      type_cast_502_inst_ack_1<= rack(0);
      type_cast_502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_556_inst_req_0;
      type_cast_556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_556_inst_req_1;
      type_cast_556_inst_ack_1<= rack(0);
      type_cast_556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_574_inst_req_0;
      type_cast_574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_574_inst_req_1;
      type_cast_574_inst_ack_1<= rack(0);
      type_cast_574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_641_inst_req_0;
      type_cast_641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_641_inst_req_1;
      type_cast_641_inst_ack_1<= rack(0);
      type_cast_641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_641_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp491x_xop_638,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_38_642,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_664_inst_req_0;
      type_cast_664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_664_inst_req_1;
      type_cast_664_inst_ack_1<= rack(0);
      type_cast_664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext483_815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_664_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_678_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_678_inst_req_0;
      type_cast_678_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_678_inst_req_1;
      type_cast_678_inst_ack_1<= rack(0);
      type_cast_678_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_678_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_691_inst_req_0;
      type_cast_691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_691_inst_req_1;
      type_cast_691_inst_ack_1<= rack(0);
      type_cast_691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_688,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_745_inst_req_0;
      type_cast_745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_745_inst_req_1;
      type_cast_745_inst_ack_1<= rack(0);
      type_cast_745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_763_inst_req_1;
      type_cast_763_inst_ack_1<= rack(0);
      type_cast_763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_832_inst_req_0;
      type_cast_832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_832_inst_req_1;
      type_cast_832_inst_ack_1<= rack(0);
      type_cast_832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_836_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_836_inst_req_0;
      type_cast_836_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_836_inst_req_1;
      type_cast_836_inst_ack_1<= rack(0);
      type_cast_836_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_836_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_837,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_840_inst_req_0;
      type_cast_840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_840_inst_req_1;
      type_cast_840_inst_ack_1<= rack(0);
      type_cast_840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_841,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_885_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_885_inst_req_0;
      type_cast_885_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_885_inst_req_1;
      type_cast_885_inst_ack_1<= rack(0);
      type_cast_885_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_885_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp475x_xop_882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_886,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_908_inst_req_0;
      type_cast_908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_908_inst_req_1;
      type_cast_908_inst_ack_1<= rack(0);
      type_cast_908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext469_927,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_908_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_949_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_949_inst_req_0;
      type_cast_949_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_949_inst_req_1;
      type_cast_949_inst_ack_1<= rack(0);
      type_cast_949_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_949_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_948_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_950,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1168_index_1_rename
    process(R_indvar_1167_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1167_resized;
      ov(13 downto 0) := iv;
      R_indvar_1167_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1168_index_1_resize
    process(indvar_1156) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1156;
      ov := iv(13 downto 0);
      R_indvar_1167_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1168_root_address_inst
    process(array_obj_ref_1168_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1168_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1168_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_index_1_rename
    process(R_indvar498_462_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar498_462_resized;
      ov(13 downto 0) := iv;
      R_indvar498_462_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_index_1_resize
    process(indvar498_451) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar498_451;
      ov := iv(13 downto 0);
      R_indvar498_462_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_root_address_inst
    process(array_obj_ref_463_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_463_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_463_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_670_index_1_rename
    process(R_indvar482_669_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar482_669_resized;
      ov(10 downto 0) := iv;
      R_indvar482_669_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_670_index_1_resize
    process(indvar482_658) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar482_658;
      ov := iv(10 downto 0);
      R_indvar482_669_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_670_root_address_inst
    process(array_obj_ref_670_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_670_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_670_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_914_index_1_rename
    process(R_indvar468_913_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar468_913_resized;
      ov(13 downto 0) := iv;
      R_indvar468_913_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_914_index_1_resize
    process(indvar468_902) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar468_902;
      ov := iv(13 downto 0);
      R_indvar468_913_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_914_root_address_inst
    process(array_obj_ref_914_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_914_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_914_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1173_addr_0
    process(ptr_deref_1173_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1173_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1173_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1173_base_resize
    process(arrayidx375_1170) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx375_1170;
      ov := iv(13 downto 0);
      ptr_deref_1173_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1173_gather_scatter
    process(ptr_deref_1173_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1173_data_0;
      ov(63 downto 0) := iv;
      tmp376_1174 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1173_root_address_inst
    process(ptr_deref_1173_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1173_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1173_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_600_addr_0
    process(ptr_deref_600_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_600_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_600_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_600_base_resize
    process(arrayidx_465) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_465;
      ov := iv(13 downto 0);
      ptr_deref_600_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_600_gather_scatter
    process(add186_598) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_598;
      ov(63 downto 0) := iv;
      ptr_deref_600_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_600_root_address_inst
    process(ptr_deref_600_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_600_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_600_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_addr_0
    process(ptr_deref_807_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_807_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_807_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_base_resize
    process(arrayidx246_672) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_672;
      ov := iv(10 downto 0);
      ptr_deref_807_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_gather_scatter
    process(add242_805) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_805;
      ov(63 downto 0) := iv;
      ptr_deref_807_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_root_address_inst
    process(ptr_deref_807_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_807_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_807_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_918_addr_0
    process(ptr_deref_918_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_918_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_918_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_918_base_resize
    process(arrayidx269_916) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_916;
      ov := iv(13 downto 0);
      ptr_deref_918_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_918_gather_scatter
    process(type_cast_920_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_920_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_918_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_918_root_address_inst
    process(ptr_deref_918_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_918_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_918_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1112_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264448_857;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1112_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1112_branch_req_0,
          ack0 => if_stmt_1112_branch_ack_0,
          ack1 => if_stmt_1112_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1284_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1283;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1284_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1284_branch_req_0,
          ack0 => if_stmt_1284_branch_ack_0,
          ack1 => if_stmt_1284_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_392_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp456_391;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_392_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_392_branch_req_0,
          ack0 => if_stmt_392_branch_ack_0,
          ack1 => if_stmt_392_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_407_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194452_406;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_407_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_407_branch_req_0,
          ack0 => if_stmt_407_branch_ack_0,
          ack1 => if_stmt_407_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_614_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_613;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_614_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_614_branch_req_0,
          ack0 => if_stmt_614_branch_ack_0,
          ack1 => if_stmt_614_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_821_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_820;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_821_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_821_branch_req_0,
          ack0 => if_stmt_821_branch_ack_0,
          ack1 => if_stmt_821_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_858_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264448_857;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_858_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_858_branch_req_0,
          ack0 => if_stmt_858_branch_ack_0,
          ack1 => if_stmt_858_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_933_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_932;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_933_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_933_branch_req_0,
          ack0 => if_stmt_933_branch_ack_0,
          ack1 => if_stmt_933_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1135_inst
    process(tmp463_1124) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp463_1124, type_cast_1134_wire_constant, tmp_var);
      tmp463x_xop_1136 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_430_inst
    process(tmp505_419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp505_419, type_cast_429_wire_constant, tmp_var);
      tmp505x_xop_431 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_637_inst
    process(tmp491_626) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp491_626, type_cast_636_wire_constant, tmp_var);
      tmp491x_xop_638 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_881_inst
    process(tmp475_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp475_870, type_cast_880_wire_constant, tmp_var);
      tmp475x_xop_882 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1145_inst
    process(iNsTr_108_1140) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_108_1140, type_cast_1144_wire_constant, tmp_var);
      xx_xop_1146 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1277_inst
    process(indvar_1156) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1156, type_cast_1276_wire_constant, tmp_var);
      indvarx_xnext_1278 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_440_inst
    process(iNsTr_25_435) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_25_435, type_cast_439_wire_constant, tmp_var);
      xx_xop514_441 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_607_inst
    process(indvar498_451) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar498_451, type_cast_606_wire_constant, tmp_var);
      indvarx_xnext499_608 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_647_inst
    process(iNsTr_38_642) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_38_642, type_cast_646_wire_constant, tmp_var);
      xx_xop513_648 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_814_inst
    process(indvar482_658) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar482_658, type_cast_813_wire_constant, tmp_var);
      indvarx_xnext483_815 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_891_inst
    process(iNsTr_52_886) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_52_886, type_cast_890_wire_constant, tmp_var);
      xx_xop512_892 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_926_inst
    process(indvar468_902) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar468_902, type_cast_925_wire_constant, tmp_var);
      indvarx_xnext469_927 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1282_inst
    process(indvarx_xnext_1278, tmp467_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1278, tmp467_1153, tmp_var);
      exitcond1_1283 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_612_inst
    process(indvarx_xnext499_608, tmp510_448) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext499_608, tmp510_448, tmp_var);
      exitcond3_613 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_819_inst
    process(indvarx_xnext483_815, tmp496_655) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext483_815, tmp496_655, tmp_var);
      exitcond2_820 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_931_inst
    process(indvarx_xnext469_927, tmp480_899) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext469_927, tmp480_899, tmp_var);
      exitcond_932 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1123_inst
    process(mul259_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_851, type_cast_1122_wire_constant, tmp_var);
      tmp463_1124 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_418_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_417_wire_constant, tmp_var);
      tmp505_419 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_625_inst
    process(mul91_260) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_260, type_cast_624_wire_constant, tmp_var);
      tmp491_626 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_869_inst
    process(mul259_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_851, type_cast_868_wire_constant, tmp_var);
      tmp475_870 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1021_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1020_wire_constant, tmp_var);
      shr307_1022 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1031_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1030_wire_constant, tmp_var);
      shr313_1032 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1041_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1040_wire_constant, tmp_var);
      shr319_1042 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1051_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1050_wire_constant, tmp_var);
      shr325_1052 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1061_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1060_wire_constant, tmp_var);
      shr331_1062 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1071_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1070_wire_constant, tmp_var);
      shr337_1072 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1081_inst
    process(sub_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1012, type_cast_1080_wire_constant, tmp_var);
      shr343_1082 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1183_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1182_wire_constant, tmp_var);
      shr383_1184 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1193_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1192_wire_constant, tmp_var);
      shr389_1194 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1203_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1202_wire_constant, tmp_var);
      shr395_1204 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1213_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1212_wire_constant, tmp_var);
      shr401_1214 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1223_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1222_wire_constant, tmp_var);
      shr407_1224 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1233_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1232_wire_constant, tmp_var);
      shr413_1234 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1243_inst
    process(tmp376_1174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1174, type_cast_1242_wire_constant, tmp_var);
      shr419_1244 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_223_inst
    process(conv63_215, conv61_211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_215, conv61_211, tmp_var);
      mul_224 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_228_inst
    process(mul_224, conv65_219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_224, conv65_219, tmp_var);
      mul66_229 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(conv84_237, conv82_233) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_237, conv82_233, tmp_var);
      mul85_250 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_254_inst
    process(mul85_250, conv87_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_250, conv87_241, tmp_var);
      mul88_255 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_259_inst
    process(mul88_255, conv90_245) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_255, conv90_245, tmp_var);
      mul91_260 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_845_inst
    process(conv255_837, conv253_833) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_837, conv253_833, tmp_var);
      mul256_846 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_850_inst
    process(mul256_846, conv258_841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_846, conv258_841, tmp_var);
      mul259_851 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_106_inst
    process(shl18_95, conv20_102) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_95, conv20_102, tmp_var);
      add21_107 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_131_inst
    process(shl27_120, conv29_127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_120, conv29_127, tmp_var);
      add30_132 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_156_inst
    process(shl36_145, conv38_152) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_145, conv38_152, tmp_var);
      add39_157 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_181_inst
    process(shl45_170, conv47_177) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_170, conv47_177, tmp_var);
      add48_182 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_206_inst
    process(shl54_195, conv56_202) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_195, conv56_202, tmp_var);
      add57_207 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_284_inst
    process(shl96_273, conv98_280) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_273, conv98_280, tmp_var);
      add99_285 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_309_inst
    process(shl105_298, conv107_305) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_298, conv107_305, tmp_var);
      add108_310 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_334_inst
    process(shl114_323, conv116_330) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_323, conv116_330, tmp_var);
      add117_335 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_359_inst
    process(shl123_348, conv125_355) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_348, conv125_355, tmp_var);
      add126_360 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_384_inst
    process(shl132_373, conv134_380) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_373, conv134_380, tmp_var);
      add135_385 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_56_inst
    process(shl_45, conv3_52) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_45, conv3_52, tmp_var);
      add_57 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_81_inst
    process(shl9_70, conv11_77) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_70, conv11_77, tmp_var);
      add12_82 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_489_inst
    process(shl146_478, conv149_485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_478, conv149_485, tmp_var);
      add150_490 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_507_inst
    process(shl152_496, conv155_503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_496, conv155_503, tmp_var);
      add156_508 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_525_inst
    process(shl158_514, conv161_521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_514, conv161_521, tmp_var);
      add162_526 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_543_inst
    process(shl164_532, conv167_539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_532, conv167_539, tmp_var);
      add168_544 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_561_inst
    process(shl170_550, conv173_557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_550, conv173_557, tmp_var);
      add174_562 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_579_inst
    process(shl176_568, conv179_575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_568, conv179_575, tmp_var);
      add180_580 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_597_inst
    process(shl182_586, conv185_593) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_586, conv185_593, tmp_var);
      add186_598 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_696_inst
    process(shl202_685, conv205_692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_685, conv205_692, tmp_var);
      add206_697 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_714_inst
    process(shl208_703, conv211_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_703, conv211_710, tmp_var);
      add212_715 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_732_inst
    process(shl214_721, conv217_728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_721, conv217_728, tmp_var);
      add218_733 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_750_inst
    process(shl220_739, conv223_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_739, conv223_746, tmp_var);
      add224_751 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_768_inst
    process(shl226_757, conv229_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_757, conv229_764, tmp_var);
      add230_769 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_786_inst
    process(shl232_775, conv235_782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_775, conv235_782, tmp_var);
      add236_787 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_804_inst
    process(shl238_793, conv241_800) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_793, conv241_800, tmp_var);
      add242_805 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_119_inst
    process(conv26_114) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_114, type_cast_118_wire_constant, tmp_var);
      shl27_120 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_144_inst
    process(conv35_139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_139, type_cast_143_wire_constant, tmp_var);
      shl36_145 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_169_inst
    process(conv44_164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_164, type_cast_168_wire_constant, tmp_var);
      shl45_170 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_194_inst
    process(conv53_189) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_189, type_cast_193_wire_constant, tmp_var);
      shl54_195 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_272_inst
    process(conv95_267) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_267, type_cast_271_wire_constant, tmp_var);
      shl96_273 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_297_inst
    process(conv104_292) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_292, type_cast_296_wire_constant, tmp_var);
      shl105_298 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_322_inst
    process(conv113_317) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_317, type_cast_321_wire_constant, tmp_var);
      shl114_323 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_347_inst
    process(conv122_342) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_342, type_cast_346_wire_constant, tmp_var);
      shl123_348 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_372_inst
    process(conv131_367) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_367, type_cast_371_wire_constant, tmp_var);
      shl132_373 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_44_inst
    process(conv1_39) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_39, type_cast_43_wire_constant, tmp_var);
      shl_45 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_69_inst
    process(conv8_64) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_64, type_cast_68_wire_constant, tmp_var);
      shl9_70 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_94_inst
    process(conv17_89) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_89, type_cast_93_wire_constant, tmp_var);
      shl18_95 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_477_inst
    process(conv144_472) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_472, type_cast_476_wire_constant, tmp_var);
      shl146_478 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_495_inst
    process(add150_490) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_490, type_cast_494_wire_constant, tmp_var);
      shl152_496 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_513_inst
    process(add156_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_508, type_cast_512_wire_constant, tmp_var);
      shl158_514 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_531_inst
    process(add162_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_526, type_cast_530_wire_constant, tmp_var);
      shl164_532 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_549_inst
    process(add168_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_544, type_cast_548_wire_constant, tmp_var);
      shl170_550 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_567_inst
    process(add174_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_562, type_cast_566_wire_constant, tmp_var);
      shl176_568 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_585_inst
    process(add180_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_580, type_cast_584_wire_constant, tmp_var);
      shl182_586 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_684_inst
    process(conv200_679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_679, type_cast_683_wire_constant, tmp_var);
      shl202_685 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_702_inst
    process(add206_697) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_697, type_cast_701_wire_constant, tmp_var);
      shl208_703 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_720_inst
    process(add212_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_715, type_cast_719_wire_constant, tmp_var);
      shl214_721 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_738_inst
    process(add218_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_733, type_cast_737_wire_constant, tmp_var);
      shl220_739 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_756_inst
    process(add224_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_751, type_cast_755_wire_constant, tmp_var);
      shl226_757 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_774_inst
    process(add230_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_769, type_cast_773_wire_constant, tmp_var);
      shl232_775 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_792_inst
    process(add236_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_787, type_cast_791_wire_constant, tmp_var);
      shl238_793 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1011_inst
    process(conv298_1007, conv276_950) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv298_1007, conv276_950, tmp_var);
      sub_1012 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1129_inst
    process(tmp463_1124) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp463_1124, type_cast_1128_wire_constant, tmp_var);
      tmp464_1130 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_390_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_229, type_cast_389_wire_constant, tmp_var);
      cmp456_391 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_405_inst
    process(mul91_260) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_260, type_cast_404_wire_constant, tmp_var);
      cmp194452_406 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_424_inst
    process(tmp505_419) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp505_419, type_cast_423_wire_constant, tmp_var);
      tmp506_425 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_631_inst
    process(tmp491_626) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp491_626, type_cast_630_wire_constant, tmp_var);
      tmp492_632 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_856_inst
    process(mul259_851) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_851, type_cast_855_wire_constant, tmp_var);
      cmp264448_857 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_875_inst
    process(tmp475_870) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp475_870, type_cast_874_wire_constant, tmp_var);
      tmp476_876 <= tmp_var; --
    end process;
    -- shared split operator group (101) : array_obj_ref_1168_index_offset 
    ApIntAdd_group_101: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1167_scaled;
      array_obj_ref_1168_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1168_index_offset_req_0;
      array_obj_ref_1168_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1168_index_offset_req_1;
      array_obj_ref_1168_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_101_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_101_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_101",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 101
    -- shared split operator group (102) : array_obj_ref_463_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar498_462_scaled;
      array_obj_ref_463_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_463_index_offset_req_0;
      array_obj_ref_463_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_463_index_offset_req_1;
      array_obj_ref_463_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : array_obj_ref_670_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar482_669_scaled;
      array_obj_ref_670_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_670_index_offset_req_0;
      array_obj_ref_670_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_670_index_offset_req_1;
      array_obj_ref_670_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : array_obj_ref_914_index_offset 
    ApIntAdd_group_104: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar468_913_scaled;
      array_obj_ref_914_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_914_index_offset_req_0;
      array_obj_ref_914_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_914_index_offset_req_1;
      array_obj_ref_914_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_104_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_104_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_104",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- unary operator type_cast_1005_inst
    process(call297_1002) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call297_1002, tmp_var);
      type_cast_1005_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_948_inst
    process(call275_944) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_944, tmp_var);
      type_cast_948_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1173_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1173_load_0_req_0;
      ptr_deref_1173_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1173_load_0_req_1;
      ptr_deref_1173_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1173_word_address_0;
      ptr_deref_1173_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_600_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_600_store_0_req_0;
      ptr_deref_600_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_600_store_0_req_1;
      ptr_deref_600_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_600_word_address_0;
      data_in <= ptr_deref_600_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_807_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_807_store_0_req_0;
      ptr_deref_807_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_807_store_0_req_1;
      ptr_deref_807_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_807_word_address_0;
      data_in <= ptr_deref_807_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(10 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_918_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_918_store_0_req_0;
      ptr_deref_918_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_918_store_0_req_1;
      ptr_deref_918_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_918_word_address_0;
      data_in <= ptr_deref_918_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_998_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_998_inst_req_0;
      RPIPE_Block0_done_998_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_998_inst_req_1;
      RPIPE_Block0_done_998_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call295_999 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_ConvTranspose_input_pipe_723_inst RPIPE_ConvTranspose_input_pipe_741_inst RPIPE_ConvTranspose_input_pipe_759_inst RPIPE_ConvTranspose_input_pipe_705_inst RPIPE_ConvTranspose_input_pipe_777_inst RPIPE_ConvTranspose_input_pipe_687_inst RPIPE_ConvTranspose_input_pipe_674_inst RPIPE_ConvTranspose_input_pipe_795_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_47_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_72_inst RPIPE_ConvTranspose_input_pipe_84_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_109_inst RPIPE_ConvTranspose_input_pipe_122_inst RPIPE_ConvTranspose_input_pipe_134_inst RPIPE_ConvTranspose_input_pipe_147_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_172_inst RPIPE_ConvTranspose_input_pipe_184_inst RPIPE_ConvTranspose_input_pipe_197_inst RPIPE_ConvTranspose_input_pipe_262_inst RPIPE_ConvTranspose_input_pipe_275_inst RPIPE_ConvTranspose_input_pipe_287_inst RPIPE_ConvTranspose_input_pipe_300_inst RPIPE_ConvTranspose_input_pipe_312_inst RPIPE_ConvTranspose_input_pipe_325_inst RPIPE_ConvTranspose_input_pipe_337_inst RPIPE_ConvTranspose_input_pipe_350_inst RPIPE_ConvTranspose_input_pipe_362_inst RPIPE_ConvTranspose_input_pipe_375_inst RPIPE_ConvTranspose_input_pipe_467_inst RPIPE_ConvTranspose_input_pipe_480_inst RPIPE_ConvTranspose_input_pipe_498_inst RPIPE_ConvTranspose_input_pipe_516_inst RPIPE_ConvTranspose_input_pipe_534_inst RPIPE_ConvTranspose_input_pipe_552_inst RPIPE_ConvTranspose_input_pipe_570_inst RPIPE_ConvTranspose_input_pipe_588_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_687_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_674_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_262_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_275_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_287_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_300_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_312_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_325_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_337_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_350_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_362_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_375_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_467_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_480_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_687_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_674_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_262_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_275_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_287_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_300_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_312_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_325_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_337_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_350_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_362_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_375_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_467_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_480_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_687_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_674_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_262_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_275_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_287_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_300_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_312_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_325_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_337_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_350_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_362_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_375_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_467_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_480_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_687_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_674_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_262_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_275_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_287_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_300_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_312_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_325_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_337_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_350_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_362_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_375_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_467_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_480_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call215_724 <= data_out(319 downto 312);
      call221_742 <= data_out(311 downto 304);
      call227_760 <= data_out(303 downto 296);
      call209_706 <= data_out(295 downto 288);
      call233_778 <= data_out(287 downto 280);
      call203_688 <= data_out(279 downto 272);
      call199_675 <= data_out(271 downto 264);
      call239_796 <= data_out(263 downto 256);
      call_35 <= data_out(255 downto 248);
      call2_48 <= data_out(247 downto 240);
      call5_60 <= data_out(239 downto 232);
      call10_73 <= data_out(231 downto 224);
      call14_85 <= data_out(223 downto 216);
      call19_98 <= data_out(215 downto 208);
      call23_110 <= data_out(207 downto 200);
      call28_123 <= data_out(199 downto 192);
      call32_135 <= data_out(191 downto 184);
      call37_148 <= data_out(183 downto 176);
      call41_160 <= data_out(175 downto 168);
      call46_173 <= data_out(167 downto 160);
      call50_185 <= data_out(159 downto 152);
      call55_198 <= data_out(151 downto 144);
      call92_263 <= data_out(143 downto 136);
      call97_276 <= data_out(135 downto 128);
      call101_288 <= data_out(127 downto 120);
      call106_301 <= data_out(119 downto 112);
      call110_313 <= data_out(111 downto 104);
      call115_326 <= data_out(103 downto 96);
      call119_338 <= data_out(95 downto 88);
      call124_351 <= data_out(87 downto 80);
      call128_363 <= data_out(79 downto 72);
      call133_376 <= data_out(71 downto 64);
      call143_468 <= data_out(63 downto 56);
      call147_481 <= data_out(55 downto 48);
      call153_499 <= data_out(47 downto 40);
      call159_517 <= data_out(39 downto 32);
      call165_535 <= data_out(31 downto 24);
      call171_553 <= data_out(23 downto 16);
      call177_571 <= data_out(15 downto 8);
      call183_589 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_1_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_1", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_Block0_start_976_inst WPIPE_Block0_start_979_inst WPIPE_Block0_start_970_inst WPIPE_Block0_start_973_inst WPIPE_Block0_start_967_inst WPIPE_Block0_start_964_inst WPIPE_Block0_start_983_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_993_inst WPIPE_Block0_start_952_inst WPIPE_Block0_start_955_inst WPIPE_Block0_start_958_inst WPIPE_Block0_start_961_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_976_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_979_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_970_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_973_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_967_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_964_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_983_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_993_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_952_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_955_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_958_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_961_inst_req_0;
      WPIPE_Block0_start_976_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_979_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_970_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_973_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_967_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_964_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_983_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_993_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_952_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_955_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_958_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_961_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_976_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_979_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_970_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_973_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_967_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_964_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_983_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_993_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_952_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_955_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_958_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_961_inst_req_1;
      WPIPE_Block0_start_976_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_979_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_970_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_973_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_967_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_964_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_983_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_993_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_952_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_955_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_958_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_961_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add108_310 & type_cast_981_wire_constant & add57_207 & add99_285 & add48_182 & add39_157 & type_cast_985_wire_constant & add117_335 & add126_360 & add135_385 & add_57 & add12_82 & add21_107 & add30_132;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_ConvTranspose_output_pipe_1108_inst WPIPE_ConvTranspose_output_pipe_1093_inst WPIPE_ConvTranspose_output_pipe_1099_inst WPIPE_ConvTranspose_output_pipe_1102_inst WPIPE_ConvTranspose_output_pipe_1105_inst WPIPE_ConvTranspose_output_pipe_1096_inst WPIPE_ConvTranspose_output_pipe_1087_inst WPIPE_ConvTranspose_output_pipe_1090_inst WPIPE_ConvTranspose_output_pipe_1249_inst WPIPE_ConvTranspose_output_pipe_1252_inst WPIPE_ConvTranspose_output_pipe_1255_inst WPIPE_ConvTranspose_output_pipe_1258_inst WPIPE_ConvTranspose_output_pipe_1261_inst WPIPE_ConvTranspose_output_pipe_1264_inst WPIPE_ConvTranspose_output_pipe_1267_inst WPIPE_ConvTranspose_output_pipe_1270_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1108_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1093_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1099_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1102_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1105_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1096_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1087_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1090_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1249_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1252_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1255_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1258_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1261_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1264_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1267_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1270_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1108_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1093_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1099_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1102_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1105_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1096_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1087_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1090_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1249_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1252_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1255_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1258_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1261_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1264_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1267_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1270_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1108_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1093_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1099_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1102_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1105_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1096_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1087_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1090_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1249_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1252_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1255_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1258_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1261_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1264_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1267_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1270_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1108_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1093_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1099_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1102_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1105_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1096_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1087_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1090_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1249_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1252_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1255_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1258_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1261_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1264_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1267_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1270_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv304_1016 & conv334_1066 & conv322_1046 & conv316_1036 & conv310_1026 & conv328_1056 & conv346_1086 & conv340_1076 & conv422_1248 & conv416_1238 & conv410_1228 & conv404_1218 & conv398_1208 & conv392_1198 & conv386_1188 & conv380_1178;
      ConvTranspose_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_1_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_944_call call_stmt_1002_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_944_call_req_0;
      reqL_unguarded(0) <= call_stmt_1002_call_req_0;
      call_stmt_944_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1002_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_944_call_req_1;
      reqR_unguarded(0) <= call_stmt_1002_call_req_1;
      call_stmt_944_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1002_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_944 <= data_out(127 downto 64);
      call297_1002 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3049_start: Boolean;
  signal convTransposeA_CP_3049_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1344_inst_req_1 : boolean;
  signal ptr_deref_1526_load_0_req_0 : boolean;
  signal ptr_deref_1526_load_0_ack_0 : boolean;
  signal RPIPE_Block0_start_1355_inst_req_0 : boolean;
  signal type_cast_1344_inst_ack_0 : boolean;
  signal type_cast_1395_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1352_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1355_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1352_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1352_inst_ack_0 : boolean;
  signal ptr_deref_1551_store_0_req_0 : boolean;
  signal ptr_deref_1551_store_0_ack_0 : boolean;
  signal type_cast_1708_inst_req_1 : boolean;
  signal type_cast_1708_inst_ack_1 : boolean;
  signal W_arrayidx72_1547_delayed_6_0_1547_inst_req_1 : boolean;
  signal W_arrayidx72_1547_delayed_6_0_1547_inst_ack_1 : boolean;
  signal W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_ack_0 : boolean;
  signal add_dest_dim0x_x1_at_entry_1419_1454_buf_req_0 : boolean;
  signal add_dest_dim0x_x1_at_entry_1419_1454_buf_ack_0 : boolean;
  signal phi_stmt_1455_req_0 : boolean;
  signal phi_stmt_1450_req_1 : boolean;
  signal add_dest_dim0x_x1_at_entry_1419_1454_buf_req_1 : boolean;
  signal RPIPE_Block0_start_1355_inst_req_1 : boolean;
  signal type_cast_1395_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1355_inst_ack_1 : boolean;
  signal phi_stmt_1450_ack_0 : boolean;
  signal phi_stmt_1455_req_1 : boolean;
  signal type_cast_1680_inst_req_0 : boolean;
  signal W_arrayidx72_1547_delayed_6_0_1547_inst_ack_0 : boolean;
  signal type_cast_1344_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1358_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1358_inst_ack_0 : boolean;
  signal type_cast_1449_inst_req_0 : boolean;
  signal type_cast_1453_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1358_inst_req_1 : boolean;
  signal phi_stmt_1455_ack_0 : boolean;
  signal RPIPE_Block0_start_1358_inst_ack_1 : boolean;
  signal W_input_dim1x_x1_1599_delayed_2_0_1609_inst_ack_1 : boolean;
  signal W_arrayidx72_1547_delayed_6_0_1547_inst_req_0 : boolean;
  signal type_cast_1453_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1340_inst_req_0 : boolean;
  signal phi_stmt_1445_req_1 : boolean;
  signal type_cast_1379_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1340_inst_ack_0 : boolean;
  signal type_cast_1449_inst_ack_0 : boolean;
  signal type_cast_1379_inst_ack_0 : boolean;
  signal type_cast_1453_inst_req_0 : boolean;
  signal type_cast_1404_inst_req_1 : boolean;
  signal type_cast_1404_inst_ack_1 : boolean;
  signal phi_stmt_1445_req_0 : boolean;
  signal type_cast_1449_inst_req_1 : boolean;
  signal type_cast_1379_inst_req_1 : boolean;
  signal type_cast_1379_inst_ack_1 : boolean;
  signal type_cast_1449_inst_ack_1 : boolean;
  signal type_cast_1453_inst_ack_0 : boolean;
  signal ptr_deref_1526_load_0_ack_1 : boolean;
  signal type_cast_1395_inst_req_0 : boolean;
  signal phi_stmt_1450_req_0 : boolean;
  signal phi_stmt_1445_ack_0 : boolean;
  signal W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_req_0 : boolean;
  signal type_cast_1458_inst_req_0 : boolean;
  signal type_cast_1458_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1340_inst_req_1 : boolean;
  signal type_cast_1395_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1352_inst_req_0 : boolean;
  signal type_cast_1383_inst_req_0 : boolean;
  signal type_cast_1383_inst_ack_0 : boolean;
  signal add_dest_dim0x_x1_at_entry_1419_1454_buf_ack_1 : boolean;
  signal type_cast_1404_inst_req_0 : boolean;
  signal type_cast_1383_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1340_inst_ack_1 : boolean;
  signal type_cast_1344_inst_req_0 : boolean;
  signal type_cast_1383_inst_ack_1 : boolean;
  signal type_cast_1404_inst_ack_0 : boolean;
  signal W_input_dim1x_x1_1599_delayed_2_0_1609_inst_req_1 : boolean;
  signal type_cast_1331_inst_ack_1 : boolean;
  signal type_cast_1331_inst_req_1 : boolean;
  signal do_while_stmt_1443_branch_req_0 : boolean;
  signal if_stmt_1742_branch_req_0 : boolean;
  signal addr_of_1522_final_reg_req_1 : boolean;
  signal ptr_deref_1526_load_0_req_1 : boolean;
  signal type_cast_1601_inst_req_0 : boolean;
  signal addr_of_1522_final_reg_ack_1 : boolean;
  signal RPIPE_Block0_start_1300_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1300_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1300_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1300_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1303_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1303_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1303_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1303_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1306_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1306_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1306_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1306_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1309_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1309_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1309_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1309_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1312_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1312_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1312_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1312_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1315_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1315_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1315_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1315_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1318_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1318_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1318_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1318_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1321_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1321_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1321_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1321_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1324_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1324_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1324_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1324_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1327_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1327_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1327_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1327_inst_ack_1 : boolean;
  signal type_cast_1331_inst_req_0 : boolean;
  signal type_cast_1331_inst_ack_0 : boolean;
  signal type_cast_1458_inst_req_1 : boolean;
  signal type_cast_1458_inst_ack_1 : boolean;
  signal type_cast_1723_inst_ack_1 : boolean;
  signal addr_of_1545_final_reg_ack_1 : boolean;
  signal addr_of_1545_final_reg_req_1 : boolean;
  signal add_dest_dim1x_x1_at_entry_1423_1459_buf_req_0 : boolean;
  signal add_dest_dim1x_x1_at_entry_1423_1459_buf_ack_0 : boolean;
  signal add_dest_dim1x_x1_at_entry_1423_1459_buf_req_1 : boolean;
  signal add_dest_dim1x_x1_at_entry_1423_1459_buf_ack_1 : boolean;
  signal addr_of_1545_final_reg_ack_0 : boolean;
  signal addr_of_1545_final_reg_req_0 : boolean;
  signal type_cast_1665_inst_ack_1 : boolean;
  signal type_cast_1665_inst_req_1 : boolean;
  signal phi_stmt_1460_req_0 : boolean;
  signal type_cast_1665_inst_ack_0 : boolean;
  signal type_cast_1665_inst_req_0 : boolean;
  signal phi_stmt_1460_req_1 : boolean;
  signal do_while_stmt_1443_branch_ack_1 : boolean;
  signal W_input_dim1x_x1_1599_delayed_2_0_1609_inst_ack_0 : boolean;
  signal type_cast_1560_inst_ack_1 : boolean;
  signal phi_stmt_1460_ack_0 : boolean;
  signal type_cast_1560_inst_req_1 : boolean;
  signal type_cast_1560_inst_ack_0 : boolean;
  signal type_cast_1560_inst_req_0 : boolean;
  signal type_cast_1463_inst_req_0 : boolean;
  signal type_cast_1463_inst_ack_0 : boolean;
  signal type_cast_1463_inst_req_1 : boolean;
  signal type_cast_1463_inst_ack_1 : boolean;
  signal type_cast_1708_inst_ack_0 : boolean;
  signal type_cast_1723_inst_req_1 : boolean;
  signal W_input_dim1x_x1_1599_delayed_2_0_1609_inst_req_0 : boolean;
  signal W_add87_1582_delayed_1_0_1589_inst_ack_1 : boolean;
  signal W_add87_1582_delayed_1_0_1589_inst_req_1 : boolean;
  signal W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_ack_1 : boolean;
  signal W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_req_1 : boolean;
  signal phi_stmt_1465_req_0 : boolean;
  signal phi_stmt_1465_req_1 : boolean;
  signal W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_ack_0 : boolean;
  signal W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_req_0 : boolean;
  signal phi_stmt_1465_ack_0 : boolean;
  signal type_cast_1556_inst_ack_1 : boolean;
  signal type_cast_1556_inst_req_1 : boolean;
  signal array_obj_ref_1544_index_offset_ack_1 : boolean;
  signal type_cast_1468_inst_req_0 : boolean;
  signal type_cast_1468_inst_ack_0 : boolean;
  signal type_cast_1468_inst_req_1 : boolean;
  signal type_cast_1468_inst_ack_1 : boolean;
  signal type_cast_1708_inst_req_0 : boolean;
  signal array_obj_ref_1544_index_offset_req_1 : boolean;
  signal W_add87_1582_delayed_1_0_1589_inst_ack_0 : boolean;
  signal W_add87_1582_delayed_1_0_1589_inst_req_0 : boolean;
  signal array_obj_ref_1544_index_offset_ack_0 : boolean;
  signal array_obj_ref_1544_index_offset_req_0 : boolean;
  signal W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_ack_1 : boolean;
  signal W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_req_1 : boolean;
  signal phi_stmt_1470_req_0 : boolean;
  signal W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_ack_0 : boolean;
  signal phi_stmt_1470_req_1 : boolean;
  signal W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_req_0 : boolean;
  signal phi_stmt_1470_ack_0 : boolean;
  signal type_cast_1556_inst_ack_0 : boolean;
  signal type_cast_1556_inst_req_0 : boolean;
  signal type_cast_1473_inst_req_0 : boolean;
  signal type_cast_1473_inst_ack_0 : boolean;
  signal type_cast_1473_inst_req_1 : boolean;
  signal type_cast_1473_inst_ack_1 : boolean;
  signal do_while_stmt_1443_branch_ack_0 : boolean;
  signal W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_ack_1 : boolean;
  signal W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_req_1 : boolean;
  signal type_cast_1680_inst_ack_1 : boolean;
  signal type_cast_1680_inst_req_1 : boolean;
  signal type_cast_1680_inst_ack_0 : boolean;
  signal type_cast_1601_inst_ack_1 : boolean;
  signal type_cast_1483_inst_req_0 : boolean;
  signal type_cast_1483_inst_ack_0 : boolean;
  signal W_input_dim0x_x1_1619_delayed_2_0_1632_inst_ack_1 : boolean;
  signal type_cast_1483_inst_req_1 : boolean;
  signal type_cast_1483_inst_ack_1 : boolean;
  signal type_cast_1723_inst_ack_0 : boolean;
  signal type_cast_1601_inst_req_1 : boolean;
  signal W_input_dim0x_x1_1619_delayed_2_0_1632_inst_req_1 : boolean;
  signal addr_of_1522_final_reg_ack_0 : boolean;
  signal type_cast_1487_inst_req_0 : boolean;
  signal type_cast_1487_inst_ack_0 : boolean;
  signal type_cast_1487_inst_req_1 : boolean;
  signal type_cast_1487_inst_ack_1 : boolean;
  signal type_cast_1723_inst_req_0 : boolean;
  signal W_input_dim0x_x1_1619_delayed_2_0_1632_inst_ack_0 : boolean;
  signal addr_of_1522_final_reg_req_0 : boolean;
  signal W_input_dim0x_x1_1619_delayed_2_0_1632_inst_req_0 : boolean;
  signal type_cast_1491_inst_req_0 : boolean;
  signal type_cast_1491_inst_ack_0 : boolean;
  signal type_cast_1491_inst_req_1 : boolean;
  signal type_cast_1491_inst_ack_1 : boolean;
  signal ptr_deref_1551_store_0_ack_1 : boolean;
  signal type_cast_1515_inst_req_0 : boolean;
  signal type_cast_1515_inst_ack_0 : boolean;
  signal type_cast_1515_inst_req_1 : boolean;
  signal type_cast_1515_inst_ack_1 : boolean;
  signal type_cast_1601_inst_ack_0 : boolean;
  signal ptr_deref_1551_store_0_req_1 : boolean;
  signal array_obj_ref_1521_index_offset_req_0 : boolean;
  signal array_obj_ref_1521_index_offset_ack_0 : boolean;
  signal array_obj_ref_1521_index_offset_req_1 : boolean;
  signal array_obj_ref_1521_index_offset_ack_1 : boolean;
  signal if_stmt_1742_branch_ack_1 : boolean;
  signal if_stmt_1742_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1748_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1748_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1748_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1748_inst_ack_1 : boolean;
  signal type_cast_1426_inst_req_0 : boolean;
  signal type_cast_1426_inst_ack_0 : boolean;
  signal type_cast_1426_inst_req_1 : boolean;
  signal type_cast_1426_inst_ack_1 : boolean;
  signal phi_stmt_1423_req_0 : boolean;
  signal type_cast_1422_inst_req_0 : boolean;
  signal type_cast_1422_inst_ack_0 : boolean;
  signal type_cast_1422_inst_req_1 : boolean;
  signal type_cast_1422_inst_ack_1 : boolean;
  signal phi_stmt_1419_req_0 : boolean;
  signal phi_stmt_1419_ack_0 : boolean;
  signal phi_stmt_1423_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3049_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3049_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3049_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3049_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3049: Block -- control-path 
    signal convTransposeA_CP_3049_elements: BooleanArray(294 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3049_elements(0) <= convTransposeA_CP_3049_start;
    convTransposeA_CP_3049_symbol <= convTransposeA_CP_3049_elements(284);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1298/$entry
      -- CP-element group 0: 	 branch_block_stmt_1298/branch_block_stmt_1298__entry__
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359__entry__
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/$entry
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_update_start_
      -- 
    cr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(0), ack => type_cast_1344_inst_req_1); -- 
    cr_3228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(0), ack => type_cast_1331_inst_req_1); -- 
    rr_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(0), ack => RPIPE_Block0_start_1300_inst_req_0); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	280 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	281 
    -- CP-element group 1: 	282 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1298/R_ifx_xend122_whilex_xend_taken_1743_place
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1298/do_while_stmt_1443__exit__
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742__entry__
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1298/if_stmt_1742_else_link/$entry
      -- 
    branch_req_4124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(1), ack => if_stmt_1742_branch_req_0); -- 
    convTransposeA_CP_3049_elements(1) <= convTransposeA_CP_3049_elements(280);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Update/cr
      -- 
    ra_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1300_inst_ack_0, ack => convTransposeA_CP_3049_elements(2)); -- 
    cr_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(2), ack => RPIPE_Block0_start_1300_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1300_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Sample/rr
      -- 
    ca_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1300_inst_ack_1, ack => convTransposeA_CP_3049_elements(3)); -- 
    rr_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(3), ack => RPIPE_Block0_start_1303_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Update/cr
      -- 
    ra_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1303_inst_ack_0, ack => convTransposeA_CP_3049_elements(4)); -- 
    cr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(4), ack => RPIPE_Block0_start_1303_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1303_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Sample/rr
      -- 
    ca_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1303_inst_ack_1, ack => convTransposeA_CP_3049_elements(5)); -- 
    rr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(5), ack => RPIPE_Block0_start_1306_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Update/cr
      -- 
    ra_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1306_inst_ack_0, ack => convTransposeA_CP_3049_elements(6)); -- 
    cr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(6), ack => RPIPE_Block0_start_1306_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1306_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Sample/rr
      -- 
    ca_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1306_inst_ack_1, ack => convTransposeA_CP_3049_elements(7)); -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(7), ack => RPIPE_Block0_start_1309_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Update/cr
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1309_inst_ack_0, ack => convTransposeA_CP_3049_elements(8)); -- 
    cr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(8), ack => RPIPE_Block0_start_1309_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1309_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Sample/rr
      -- 
    ca_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1309_inst_ack_1, ack => convTransposeA_CP_3049_elements(9)); -- 
    rr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(9), ack => RPIPE_Block0_start_1312_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Update/cr
      -- 
    ra_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1312_inst_ack_0, ack => convTransposeA_CP_3049_elements(10)); -- 
    cr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(10), ack => RPIPE_Block0_start_1312_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1312_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Sample/rr
      -- 
    ca_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1312_inst_ack_1, ack => convTransposeA_CP_3049_elements(11)); -- 
    rr_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(11), ack => RPIPE_Block0_start_1315_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Update/cr
      -- 
    ra_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1315_inst_ack_0, ack => convTransposeA_CP_3049_elements(12)); -- 
    cr_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(12), ack => RPIPE_Block0_start_1315_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1315_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Sample/rr
      -- 
    ca_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1315_inst_ack_1, ack => convTransposeA_CP_3049_elements(13)); -- 
    rr_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(13), ack => RPIPE_Block0_start_1318_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Update/cr
      -- 
    ra_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1318_inst_ack_0, ack => convTransposeA_CP_3049_elements(14)); -- 
    cr_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(14), ack => RPIPE_Block0_start_1318_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1318_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Sample/rr
      -- 
    ca_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1318_inst_ack_1, ack => convTransposeA_CP_3049_elements(15)); -- 
    rr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(15), ack => RPIPE_Block0_start_1321_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Update/cr
      -- 
    ra_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1321_inst_ack_0, ack => convTransposeA_CP_3049_elements(16)); -- 
    cr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(16), ack => RPIPE_Block0_start_1321_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1321_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Sample/rr
      -- 
    ca_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1321_inst_ack_1, ack => convTransposeA_CP_3049_elements(17)); -- 
    rr_3195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(17), ack => RPIPE_Block0_start_1324_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Update/cr
      -- 
    ra_3196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1324_inst_ack_0, ack => convTransposeA_CP_3049_elements(18)); -- 
    cr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(18), ack => RPIPE_Block0_start_1324_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1324_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Sample/rr
      -- 
    ca_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1324_inst_ack_1, ack => convTransposeA_CP_3049_elements(19)); -- 
    rr_3209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(19), ack => RPIPE_Block0_start_1327_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Update/cr
      -- 
    ra_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1327_inst_ack_0, ack => convTransposeA_CP_3049_elements(20)); -- 
    cr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(20), ack => RPIPE_Block0_start_1327_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1327_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Sample/rr
      -- 
    ca_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1327_inst_ack_1, ack => convTransposeA_CP_3049_elements(21)); -- 
    rr_3223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(21), ack => type_cast_1331_inst_req_0); -- 
    rr_3237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(21), ack => RPIPE_Block0_start_1340_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Sample/ra
      -- 
    ra_3224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1331_inst_ack_0, ack => convTransposeA_CP_3049_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1331_update_completed_
      -- 
    ca_3229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1331_inst_ack_1, ack => convTransposeA_CP_3049_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_sample_completed_
      -- 
    ra_3238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1340_inst_ack_0, ack => convTransposeA_CP_3049_elements(24)); -- 
    cr_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(24), ack => RPIPE_Block0_start_1340_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1340_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Sample/rr
      -- 
    ca_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1340_inst_ack_1, ack => convTransposeA_CP_3049_elements(25)); -- 
    rr_3251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(25), ack => type_cast_1344_inst_req_0); -- 
    rr_3265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(25), ack => RPIPE_Block0_start_1352_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Sample/$exit
      -- 
    ra_3252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1344_inst_ack_0, ack => convTransposeA_CP_3049_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/type_cast_1344_update_completed_
      -- 
    ca_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1344_inst_ack_1, ack => convTransposeA_CP_3049_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_update_start_
      -- 
    ra_3266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1352_inst_ack_0, ack => convTransposeA_CP_3049_elements(28)); -- 
    cr_3270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(28), ack => RPIPE_Block0_start_1352_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1352_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Sample/$entry
      -- 
    ca_3271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1352_inst_ack_1, ack => convTransposeA_CP_3049_elements(29)); -- 
    rr_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(29), ack => RPIPE_Block0_start_1355_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Update/cr
      -- 
    ra_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1355_inst_ack_0, ack => convTransposeA_CP_3049_elements(30)); -- 
    cr_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(30), ack => RPIPE_Block0_start_1355_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1355_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Sample/rr
      -- 
    ca_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1355_inst_ack_1, ack => convTransposeA_CP_3049_elements(31)); -- 
    rr_3293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(31), ack => RPIPE_Block0_start_1358_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Update/cr
      -- 
    ra_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1358_inst_ack_0, ack => convTransposeA_CP_3049_elements(32)); -- 
    cr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(32), ack => RPIPE_Block0_start_1358_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/RPIPE_Block0_start_1358_Update/ca
      -- 
    ca_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1358_inst_ack_1, ack => convTransposeA_CP_3049_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359__exit__
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411__entry__
      -- CP-element group 34: 	 branch_block_stmt_1298/assign_stmt_1301_to_assign_stmt_1359/$exit
      -- 
    cr_3343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1395_inst_req_1); -- 
    rr_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1379_inst_req_0); -- 
    cr_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1404_inst_req_1); -- 
    cr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1379_inst_req_1); -- 
    rr_3338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1395_inst_req_0); -- 
    rr_3324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1383_inst_req_0); -- 
    rr_3352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1404_inst_req_0); -- 
    cr_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(34), ack => type_cast_1383_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(23) & convTransposeA_CP_3049_elements(27) & convTransposeA_CP_3049_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_sample_completed_
      -- 
    ra_3311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_0, ack => convTransposeA_CP_3049_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1379_Update/ca
      -- 
    ca_3316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_1, ack => convTransposeA_CP_3049_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Sample/ra
      -- 
    ra_3325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1383_inst_ack_0, ack => convTransposeA_CP_3049_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1383_Update/ca
      -- 
    ca_3330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1383_inst_ack_1, ack => convTransposeA_CP_3049_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Sample/ra
      -- 
    ra_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_0, ack => convTransposeA_CP_3049_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1395_Update/$exit
      -- 
    ca_3344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_1, ack => convTransposeA_CP_3049_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Sample/ra
      -- 
    ra_3353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_0, ack => convTransposeA_CP_3049_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/type_cast_1404_Update/ca
      -- 
    ca_3358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_1, ack => convTransposeA_CP_3049_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	285 
    -- CP-element group 43: 	286 
    -- CP-element group 43: 	288 
    -- CP-element group 43: 	289 
    -- CP-element group 43:  members (20) 
      -- CP-element group 43: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411/$exit
      -- CP-element group 43: 	 branch_block_stmt_1298/assign_stmt_1366_to_assign_stmt_1411__exit__
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Update/cr
      -- 
    rr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(43), ack => type_cast_1426_inst_req_0); -- 
    cr_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(43), ack => type_cast_1426_inst_req_1); -- 
    rr_4193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(43), ack => type_cast_1422_inst_req_0); -- 
    cr_4198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(43), ack => type_cast_1422_inst_req_1); -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(36) & convTransposeA_CP_3049_elements(38) & convTransposeA_CP_3049_elements(40) & convTransposeA_CP_3049_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	294 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443__entry__
      -- CP-element group 44: 	 branch_block_stmt_1298/do_while_stmt_1443/$entry
      -- 
    convTransposeA_CP_3049_elements(44) <= convTransposeA_CP_3049_elements(294);
    -- CP-element group 45:  merge  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	280 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443__exit__
      -- 
    -- Element group convTransposeA_CP_3049_elements(45) is bound as output of CP function.
    -- CP-element group 46:  merge  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_back
      -- 
    -- Element group convTransposeA_CP_3049_elements(46) is bound as output of CP function.
    -- CP-element group 47:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	52 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	278 
    -- CP-element group 47: 	279 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1298/do_while_stmt_1443/condition_done
      -- CP-element group 47: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_taken/$entry
      -- CP-element group 47: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_exit/$entry
      -- 
    convTransposeA_CP_3049_elements(47) <= convTransposeA_CP_3049_elements(52);
    -- CP-element group 48:  branch  place  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	277 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_body_done
      -- 
    convTransposeA_CP_3049_elements(48) <= convTransposeA_CP_3049_elements(277);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	61 
    -- CP-element group 49: 	82 
    -- CP-element group 49: 	103 
    -- CP-element group 49: 	124 
    -- CP-element group 49: 	145 
    -- CP-element group 49: 	166 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/back_edge_to_loop_body
      -- 
    convTransposeA_CP_3049_elements(49) <= convTransposeA_CP_3049_elements(46);
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	44 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	63 
    -- CP-element group 50: 	84 
    -- CP-element group 50: 	105 
    -- CP-element group 50: 	126 
    -- CP-element group 50: 	147 
    -- CP-element group 50: 	168 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/first_time_through_loop_body
      -- 
    convTransposeA_CP_3049_elements(50) <= convTransposeA_CP_3049_elements(44);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	57 
    -- CP-element group 51: 	58 
    -- CP-element group 51: 	76 
    -- CP-element group 51: 	77 
    -- CP-element group 51: 	97 
    -- CP-element group 51: 	98 
    -- CP-element group 51: 	118 
    -- CP-element group 51: 	119 
    -- CP-element group 51: 	139 
    -- CP-element group 51: 	140 
    -- CP-element group 51: 	160 
    -- CP-element group 51: 	161 
    -- CP-element group 51: 	198 
    -- CP-element group 51: 	199 
    -- CP-element group 51: 	209 
    -- CP-element group 51: 	211 
    -- CP-element group 51: 	228 
    -- CP-element group 51: 	276 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/$entry
      -- CP-element group 51: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/loop_body_start
      -- 
    -- Element group convTransposeA_CP_3049_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	275 
    -- CP-element group 52: 	276 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	47 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/condition_evaluated
      -- 
    condition_evaluated_3373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(52), ack => do_while_stmt_1443_branch_req_0); -- 
    convTransposeA_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(56) & convTransposeA_CP_3049_elements(275) & convTransposeA_CP_3049_elements(276);
      gj_convTransposeA_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	57 
    -- CP-element group 53: 	76 
    -- CP-element group 53: 	97 
    -- CP-element group 53: 	118 
    -- CP-element group 53: 	139 
    -- CP-element group 53: 	160 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53: 	99 
    -- CP-element group 53: 	120 
    -- CP-element group 53: 	141 
    -- CP-element group 53: 	162 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/aggregated_phi_sample_req
      -- 
    convTransposeA_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(57) & convTransposeA_CP_3049_elements(76) & convTransposeA_CP_3049_elements(97) & convTransposeA_CP_3049_elements(118) & convTransposeA_CP_3049_elements(139) & convTransposeA_CP_3049_elements(160) & convTransposeA_CP_3049_elements(56);
      gj_convTransposeA_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	59 
    -- CP-element group 54: 	79 
    -- CP-element group 54: 	100 
    -- CP-element group 54: 	121 
    -- CP-element group 54: 	142 
    -- CP-element group 54: 	163 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	225 
    -- CP-element group 54: 	229 
    -- CP-element group 54: 	237 
    -- CP-element group 54: 	241 
    -- CP-element group 54: 	245 
    -- CP-element group 54: 	249 
    -- CP-element group 54: 	253 
    -- CP-element group 54: 	257 
    -- CP-element group 54: 	261 
    -- CP-element group 54: 	265 
    -- CP-element group 54: 	269 
    -- CP-element group 54: 	277 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: 	76 
    -- CP-element group 54: 	97 
    -- CP-element group 54: 	118 
    -- CP-element group 54: 	139 
    -- CP-element group 54: 	160 
    -- CP-element group 54:  members (7) 
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/aggregated_phi_sample_ack
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_sample_completed_
      -- 
    convTransposeA_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(59) & convTransposeA_CP_3049_elements(79) & convTransposeA_CP_3049_elements(100) & convTransposeA_CP_3049_elements(121) & convTransposeA_CP_3049_elements(142) & convTransposeA_CP_3049_elements(163);
      gj_convTransposeA_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	77 
    -- CP-element group 55: 	98 
    -- CP-element group 55: 	119 
    -- CP-element group 55: 	140 
    -- CP-element group 55: 	161 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	80 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	122 
    -- CP-element group 55: 	143 
    -- CP-element group 55: 	164 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_update_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/aggregated_phi_update_req
      -- 
    convTransposeA_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(58) & convTransposeA_CP_3049_elements(77) & convTransposeA_CP_3049_elements(98) & convTransposeA_CP_3049_elements(119) & convTransposeA_CP_3049_elements(140) & convTransposeA_CP_3049_elements(161);
      gj_convTransposeA_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	81 
    -- CP-element group 56: 	102 
    -- CP-element group 56: 	123 
    -- CP-element group 56: 	144 
    -- CP-element group 56: 	165 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/aggregated_phi_update_ack
      -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(60) & convTransposeA_CP_3049_elements(81) & convTransposeA_CP_3049_elements(102) & convTransposeA_CP_3049_elements(123) & convTransposeA_CP_3049_elements(144) & convTransposeA_CP_3049_elements(165);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	53 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_sample_start_
      -- 
    convTransposeA_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(54);
      gj_convTransposeA_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	195 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	55 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_update_start_
      -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(60) & convTransposeA_CP_3049_elements(195);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: 	193 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_update_completed__ps
      -- CP-element group 60: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_update_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	49 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_loopback_trigger
      -- 
    convTransposeA_CP_3049_elements(61) <= convTransposeA_CP_3049_elements(49);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_loopback_sample_req_ps
      -- 
    phi_stmt_1445_loopback_sample_req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1445_loopback_sample_req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(62), ack => phi_stmt_1445_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	50 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_entry_trigger
      -- 
    convTransposeA_CP_3049_elements(63) <= convTransposeA_CP_3049_elements(50);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_entry_sample_req_ps
      -- 
    phi_stmt_1445_entry_sample_req_3391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1445_entry_sample_req_3391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(64), ack => phi_stmt_1445_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1445_phi_mux_ack_ps
      -- 
    phi_stmt_1445_phi_mux_ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1445_ack_0, ack => convTransposeA_CP_3049_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_update_start_
      -- 
    -- Element group convTransposeA_CP_3049_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_update_completed__ps
      -- 
    convTransposeA_CP_3049_elements(68) <= convTransposeA_CP_3049_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_indvar_at_entry_1447_update_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_3049_elements(67), ack => convTransposeA_CP_3049_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Sample/rr
      -- 
    rr_3415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(72), ack => type_cast_1449_inst_req_0); -- 
    convTransposeA_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(70) & convTransposeA_CP_3049_elements(74);
      gj_convTransposeA_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Update/cr
      -- 
    cr_3420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(73), ack => type_cast_1449_inst_req_1); -- 
    convTransposeA_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(71) & convTransposeA_CP_3049_elements(75);
      gj_convTransposeA_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Sample/ra
      -- 
    ra_3416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1449_inst_ack_0, ack => convTransposeA_CP_3049_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1449_Update/ca
      -- 
    ca_3421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1449_inst_ack_1, ack => convTransposeA_CP_3049_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	51 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	54 
    -- CP-element group 76: 	243 
    -- CP-element group 76: 	247 
    -- CP-element group 76: 	255 
    -- CP-element group 76: 	263 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	53 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_sample_start_
      -- 
    convTransposeA_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(243) & convTransposeA_CP_3049_elements(247) & convTransposeA_CP_3049_elements(255) & convTransposeA_CP_3049_elements(263);
      gj_convTransposeA_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	51 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: 	191 
    -- CP-element group 77: 	254 
    -- CP-element group 77: 	262 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	55 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_update_start_
      -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(81) & convTransposeA_CP_3049_elements(191) & convTransposeA_CP_3049_elements(254) & convTransposeA_CP_3049_elements(262);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	53 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_sample_start__ps
      -- 
    convTransposeA_CP_3049_elements(78) <= convTransposeA_CP_3049_elements(53);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	54 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	55 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_update_start__ps
      -- 
    convTransposeA_CP_3049_elements(80) <= convTransposeA_CP_3049_elements(55);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	56 
    -- CP-element group 81: 	189 
    -- CP-element group 81: 	252 
    -- CP-element group 81: 	260 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_update_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_update_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	49 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_loopback_trigger
      -- 
    convTransposeA_CP_3049_elements(82) <= convTransposeA_CP_3049_elements(49);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_loopback_sample_req_ps
      -- 
    phi_stmt_1450_loopback_sample_req_3432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1450_loopback_sample_req_3432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(83), ack => phi_stmt_1450_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	50 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_entry_trigger
      -- 
    convTransposeA_CP_3049_elements(84) <= convTransposeA_CP_3049_elements(50);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_entry_sample_req_ps
      -- 
    phi_stmt_1450_entry_sample_req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1450_entry_sample_req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(85), ack => phi_stmt_1450_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_phi_mux_ack
      -- CP-element group 86: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1450_phi_mux_ack_ps
      -- 
    phi_stmt_1450_phi_mux_ack_3438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1450_ack_0, ack => convTransposeA_CP_3049_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_sample_start_
      -- 
    rr_3451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(89), ack => type_cast_1453_inst_req_0); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(87) & convTransposeA_CP_3049_elements(91);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_update_start_
      -- 
    cr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(90), ack => type_cast_1453_inst_req_1); -- 
    convTransposeA_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(88) & convTransposeA_CP_3049_elements(92);
      gj_convTransposeA_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Sample/ra
      -- 
    ra_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1453_inst_ack_0, ack => convTransposeA_CP_3049_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1453_update_completed_
      -- 
    ca_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1453_inst_ack_1, ack => convTransposeA_CP_3049_elements(92)); -- 
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Sample/req
      -- CP-element group 93: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Sample/$entry
      -- 
    req_3469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(93), ack => add_dest_dim0x_x1_at_entry_1419_1454_buf_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_update_start__ps
      -- 
    req_3474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(94), ack => add_dest_dim0x_x1_at_entry_1419_1454_buf_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Sample/ack
      -- CP-element group 95: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_sample_completed_
      -- 
    ack_3470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0x_x1_at_entry_1419_1454_buf_ack_0, ack => convTransposeA_CP_3049_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim0x_x1_at_entry_1454_Update/ack
      -- 
    ack_3475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0x_x1_at_entry_1419_1454_buf_ack_1, ack => convTransposeA_CP_3049_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	51 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	54 
    -- CP-element group 97: 	243 
    -- CP-element group 97: 	247 
    -- CP-element group 97: 	259 
    -- CP-element group 97: 	267 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	53 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_sample_start_
      -- 
    convTransposeA_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(243) & convTransposeA_CP_3049_elements(247) & convTransposeA_CP_3049_elements(259) & convTransposeA_CP_3049_elements(267);
      gj_convTransposeA_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	51 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: 	187 
    -- CP-element group 98: 	234 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	55 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_update_start_
      -- 
    convTransposeA_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(102) & convTransposeA_CP_3049_elements(187) & convTransposeA_CP_3049_elements(234);
      gj_convTransposeA_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	53 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_sample_start__ps
      -- 
    convTransposeA_CP_3049_elements(99) <= convTransposeA_CP_3049_elements(53);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	54 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_update_start__ps
      -- 
    convTransposeA_CP_3049_elements(101) <= convTransposeA_CP_3049_elements(55);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	56 
    -- CP-element group 102: 	185 
    -- CP-element group 102: 	232 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	49 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_loopback_trigger
      -- 
    convTransposeA_CP_3049_elements(103) <= convTransposeA_CP_3049_elements(49);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_loopback_sample_req_ps
      -- 
    phi_stmt_1455_loopback_sample_req_3486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1455_loopback_sample_req_3486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(104), ack => phi_stmt_1455_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	50 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_entry_trigger
      -- 
    convTransposeA_CP_3049_elements(105) <= convTransposeA_CP_3049_elements(50);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_entry_sample_req_ps
      -- 
    phi_stmt_1455_entry_sample_req_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1455_entry_sample_req_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(106), ack => phi_stmt_1455_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1455_phi_mux_ack_ps
      -- 
    phi_stmt_1455_phi_mux_ack_3492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1455_ack_0, ack => convTransposeA_CP_3049_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_sample_start_
      -- 
    rr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(110), ack => type_cast_1458_inst_req_0); -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(108) & convTransposeA_CP_3049_elements(112);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Update/cr
      -- 
    cr_3510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(111), ack => type_cast_1458_inst_req_1); -- 
    convTransposeA_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(109) & convTransposeA_CP_3049_elements(113);
      gj_convTransposeA_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_sample_completed_
      -- 
    ra_3506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_0, ack => convTransposeA_CP_3049_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1458_Update/ca
      -- 
    ca_3511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_1, ack => convTransposeA_CP_3049_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Sample/req
      -- 
    req_3523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(114), ack => add_dest_dim1x_x1_at_entry_1423_1459_buf_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Update/req
      -- 
    req_3528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(115), ack => add_dest_dim1x_x1_at_entry_1423_1459_buf_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Sample/ack
      -- 
    ack_3524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1x_x1_at_entry_1423_1459_buf_ack_0, ack => convTransposeA_CP_3049_elements(116)); -- 
    -- CP-element group 117:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_update_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_add_dest_dim1x_x1_at_entry_1459_Update/ack
      -- 
    ack_3529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1x_x1_at_entry_1423_1459_buf_ack_1, ack => convTransposeA_CP_3049_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	51 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	54 
    -- CP-element group 118: 	227 
    -- CP-element group 118: 	231 
    -- CP-element group 118: 	239 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	53 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_sample_start_
      -- 
    convTransposeA_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(227) & convTransposeA_CP_3049_elements(231) & convTransposeA_CP_3049_elements(239);
      gj_convTransposeA_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	51 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	183 
    -- CP-element group 119: 	226 
    -- CP-element group 119: 	238 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	55 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_update_start_
      -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(123) & convTransposeA_CP_3049_elements(183) & convTransposeA_CP_3049_elements(226) & convTransposeA_CP_3049_elements(238);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	53 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_sample_start__ps
      -- 
    convTransposeA_CP_3049_elements(120) <= convTransposeA_CP_3049_elements(53);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	54 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	55 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_update_start__ps
      -- 
    convTransposeA_CP_3049_elements(122) <= convTransposeA_CP_3049_elements(55);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	56 
    -- CP-element group 123: 	181 
    -- CP-element group 123: 	224 
    -- CP-element group 123: 	236 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	119 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	49 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_loopback_trigger
      -- 
    convTransposeA_CP_3049_elements(124) <= convTransposeA_CP_3049_elements(49);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_loopback_sample_req
      -- CP-element group 125: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_loopback_sample_req_ps
      -- 
    phi_stmt_1460_loopback_sample_req_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1460_loopback_sample_req_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(125), ack => phi_stmt_1460_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	50 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_entry_trigger
      -- 
    convTransposeA_CP_3049_elements(126) <= convTransposeA_CP_3049_elements(50);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_entry_sample_req_ps
      -- 
    phi_stmt_1460_entry_sample_req_3543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1460_entry_sample_req_3543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(127), ack => phi_stmt_1460_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1460_phi_mux_ack_ps
      -- 
    phi_stmt_1460_phi_mux_ack_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1460_ack_0, ack => convTransposeA_CP_3049_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Sample/rr
      -- 
    rr_3559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(131), ack => type_cast_1463_inst_req_0); -- 
    convTransposeA_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(129) & convTransposeA_CP_3049_elements(133);
      gj_convTransposeA_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_update_start_
      -- CP-element group 132: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Update/cr
      -- 
    cr_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(132), ack => type_cast_1463_inst_req_1); -- 
    convTransposeA_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(130) & convTransposeA_CP_3049_elements(134);
      gj_convTransposeA_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Sample/ra
      -- 
    ra_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_0, ack => convTransposeA_CP_3049_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1463_Update/ca
      -- 
    ca_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_1, ack => convTransposeA_CP_3049_elements(134)); -- 
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_sample_start__ps
      -- CP-element group 135: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_update_start__ps
      -- CP-element group 136: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_update_start_
      -- 
    -- Element group convTransposeA_CP_3049_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_update_completed__ps
      -- 
    convTransposeA_CP_3049_elements(137) <= convTransposeA_CP_3049_elements(138);
    -- CP-element group 138:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	137 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim2x_x1_at_entry_1464_update_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(138) is a control-delay.
    cp_element_138_delay: control_delay_element  generic map(name => " 138_delay", delay_value => 1)  port map(req => convTransposeA_CP_3049_elements(136), ack => convTransposeA_CP_3049_elements(138), clk => clk, reset =>reset);
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	51 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	54 
    -- CP-element group 139: 	243 
    -- CP-element group 139: 	247 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	53 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_sample_start_
      -- 
    convTransposeA_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(243) & convTransposeA_CP_3049_elements(247);
      gj_convTransposeA_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	51 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	144 
    -- CP-element group 140: 	246 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	55 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_update_start_
      -- 
    convTransposeA_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(144) & convTransposeA_CP_3049_elements(246);
      gj_convTransposeA_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	53 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_sample_start__ps
      -- 
    convTransposeA_CP_3049_elements(141) <= convTransposeA_CP_3049_elements(53);
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	54 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	55 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_update_start__ps
      -- 
    convTransposeA_CP_3049_elements(143) <= convTransposeA_CP_3049_elements(55);
    -- CP-element group 144:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	56 
    -- CP-element group 144: 	244 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	140 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	49 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_loopback_trigger
      -- 
    convTransposeA_CP_3049_elements(145) <= convTransposeA_CP_3049_elements(49);
    -- CP-element group 146:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_loopback_sample_req
      -- CP-element group 146: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_loopback_sample_req_ps
      -- 
    phi_stmt_1465_loopback_sample_req_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1465_loopback_sample_req_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(146), ack => phi_stmt_1465_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(146) is bound as output of CP function.
    -- CP-element group 147:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	50 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_entry_trigger
      -- 
    convTransposeA_CP_3049_elements(147) <= convTransposeA_CP_3049_elements(50);
    -- CP-element group 148:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_entry_sample_req
      -- CP-element group 148: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_entry_sample_req_ps
      -- 
    phi_stmt_1465_entry_sample_req_3587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1465_entry_sample_req_3587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(148), ack => phi_stmt_1465_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_phi_mux_ack
      -- CP-element group 149: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1465_phi_mux_ack_ps
      -- 
    phi_stmt_1465_phi_mux_ack_3590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1465_ack_0, ack => convTransposeA_CP_3049_elements(149)); -- 
    -- CP-element group 150:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Sample/rr
      -- 
    rr_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(152), ack => type_cast_1468_inst_req_0); -- 
    convTransposeA_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(150) & convTransposeA_CP_3049_elements(154);
      gj_convTransposeA_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_update_start_
      -- CP-element group 153: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Update/cr
      -- 
    cr_3608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(153), ack => type_cast_1468_inst_req_1); -- 
    convTransposeA_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(151) & convTransposeA_CP_3049_elements(155);
      gj_convTransposeA_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_sample_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Sample/ra
      -- 
    ra_3604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_0, ack => convTransposeA_CP_3049_elements(154)); -- 
    -- CP-element group 155:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_update_completed__ps
      -- CP-element group 155: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1468_Update/ca
      -- 
    ca_3609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_1, ack => convTransposeA_CP_3049_elements(155)); -- 
    -- CP-element group 156:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (4) 
      -- CP-element group 156: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_sample_start__ps
      -- CP-element group 156: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_sample_completed__ps
      -- CP-element group 156: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(156) is bound as output of CP function.
    -- CP-element group 157:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (2) 
      -- CP-element group 157: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_update_start__ps
      -- CP-element group 157: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_update_start_
      -- 
    -- Element group convTransposeA_CP_3049_elements(157) is bound as output of CP function.
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_update_completed__ps
      -- 
    convTransposeA_CP_3049_elements(158) <= convTransposeA_CP_3049_elements(159);
    -- CP-element group 159:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	158 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim1x_x1_at_entry_1469_update_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(159) is a control-delay.
    cp_element_159_delay: control_delay_element  generic map(name => " 159_delay", delay_value => 1)  port map(req => convTransposeA_CP_3049_elements(157), ack => convTransposeA_CP_3049_elements(159), clk => clk, reset =>reset);
    -- CP-element group 160:  join  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	51 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	54 
    -- CP-element group 160: 	243 
    -- CP-element group 160: 	247 
    -- CP-element group 160: 	251 
    -- CP-element group 160: 	271 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	53 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_sample_start_
      -- 
    convTransposeA_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(243) & convTransposeA_CP_3049_elements(247) & convTransposeA_CP_3049_elements(251) & convTransposeA_CP_3049_elements(271);
      gj_convTransposeA_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	51 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	165 
    -- CP-element group 161: 	250 
    -- CP-element group 161: 	270 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	55 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_update_start_
      -- 
    convTransposeA_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(165) & convTransposeA_CP_3049_elements(250) & convTransposeA_CP_3049_elements(270);
      gj_convTransposeA_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	53 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_sample_start__ps
      -- 
    convTransposeA_CP_3049_elements(162) <= convTransposeA_CP_3049_elements(53);
    -- CP-element group 163:  join  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	54 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(163) is bound as output of CP function.
    -- CP-element group 164:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	55 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_update_start__ps
      -- 
    convTransposeA_CP_3049_elements(164) <= convTransposeA_CP_3049_elements(55);
    -- CP-element group 165:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	56 
    -- CP-element group 165: 	248 
    -- CP-element group 165: 	268 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	161 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(165) is bound as output of CP function.
    -- CP-element group 166:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	49 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_loopback_trigger
      -- 
    convTransposeA_CP_3049_elements(166) <= convTransposeA_CP_3049_elements(49);
    -- CP-element group 167:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_loopback_sample_req
      -- CP-element group 167: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_loopback_sample_req_ps
      -- 
    phi_stmt_1470_loopback_sample_req_3628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1470_loopback_sample_req_3628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(167), ack => phi_stmt_1470_req_0); -- 
    -- Element group convTransposeA_CP_3049_elements(167) is bound as output of CP function.
    -- CP-element group 168:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	50 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_entry_trigger
      -- 
    convTransposeA_CP_3049_elements(168) <= convTransposeA_CP_3049_elements(50);
    -- CP-element group 169:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_entry_sample_req
      -- CP-element group 169: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_entry_sample_req_ps
      -- 
    phi_stmt_1470_entry_sample_req_3631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1470_entry_sample_req_3631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(169), ack => phi_stmt_1470_req_1); -- 
    -- Element group convTransposeA_CP_3049_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_phi_mux_ack
      -- CP-element group 170: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/phi_stmt_1470_phi_mux_ack_ps
      -- 
    phi_stmt_1470_phi_mux_ack_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1470_ack_0, ack => convTransposeA_CP_3049_elements(170)); -- 
    -- CP-element group 171:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (1) 
      -- CP-element group 172: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3049_elements(172) is bound as output of CP function.
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Sample/rr
      -- 
    rr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(173), ack => type_cast_1473_inst_req_0); -- 
    convTransposeA_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(171) & convTransposeA_CP_3049_elements(175);
      gj_convTransposeA_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_update_start_
      -- CP-element group 174: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Update/cr
      -- 
    cr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(174), ack => type_cast_1473_inst_req_1); -- 
    convTransposeA_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(172) & convTransposeA_CP_3049_elements(176);
      gj_convTransposeA_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (4) 
      -- CP-element group 175: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_sample_completed__ps
      -- CP-element group 175: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Sample/ra
      -- 
    ra_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1473_inst_ack_0, ack => convTransposeA_CP_3049_elements(175)); -- 
    -- CP-element group 176:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (4) 
      -- CP-element group 176: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_update_completed__ps
      -- CP-element group 176: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1473_Update/ca
      -- 
    ca_3653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1473_inst_ack_1, ack => convTransposeA_CP_3049_elements(176)); -- 
    -- CP-element group 177:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (4) 
      -- CP-element group 177: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_sample_start__ps
      -- CP-element group 177: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_sample_completed__ps
      -- CP-element group 177: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(177) is bound as output of CP function.
    -- CP-element group 178:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_update_start__ps
      -- CP-element group 178: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_update_start_
      -- 
    -- Element group convTransposeA_CP_3049_elements(178) is bound as output of CP function.
    -- CP-element group 179:  join  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_update_completed__ps
      -- 
    convTransposeA_CP_3049_elements(179) <= convTransposeA_CP_3049_elements(180);
    -- CP-element group 180:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	179 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/R_input_dim0x_x1_at_entry_1474_update_completed_
      -- 
    -- Element group convTransposeA_CP_3049_elements(180) is a control-delay.
    cp_element_180_delay: control_delay_element  generic map(name => " 180_delay", delay_value => 1)  port map(req => convTransposeA_CP_3049_elements(178), ack => convTransposeA_CP_3049_elements(180), clk => clk, reset =>reset);
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	123 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Sample/rr
      -- 
    rr_3670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(181), ack => type_cast_1483_inst_req_0); -- 
    convTransposeA_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(123) & convTransposeA_CP_3049_elements(183);
      gj_convTransposeA_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	212 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_update_start_
      -- CP-element group 182: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Update/cr
      -- 
    cr_3675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(182), ack => type_cast_1483_inst_req_1); -- 
    convTransposeA_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(184) & convTransposeA_CP_3049_elements(212);
      gj_convTransposeA_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	119 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Sample/ra
      -- 
    ra_3671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1483_inst_ack_0, ack => convTransposeA_CP_3049_elements(183)); -- 
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	210 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1483_Update/ca
      -- 
    ca_3676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1483_inst_ack_1, ack => convTransposeA_CP_3049_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	102 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Sample/rr
      -- 
    rr_3684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(185), ack => type_cast_1487_inst_req_0); -- 
    convTransposeA_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(102) & convTransposeA_CP_3049_elements(187);
      gj_convTransposeA_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: 	212 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_update_start_
      -- CP-element group 186: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Update/cr
      -- 
    cr_3689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(186), ack => type_cast_1487_inst_req_1); -- 
    convTransposeA_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(188) & convTransposeA_CP_3049_elements(212);
      gj_convTransposeA_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	98 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Sample/ra
      -- 
    ra_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1487_inst_ack_0, ack => convTransposeA_CP_3049_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	210 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1487_Update/ca
      -- 
    ca_3690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1487_inst_ack_1, ack => convTransposeA_CP_3049_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	81 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Sample/rr
      -- 
    rr_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(189), ack => type_cast_1491_inst_req_0); -- 
    convTransposeA_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(81) & convTransposeA_CP_3049_elements(191);
      gj_convTransposeA_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	212 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_update_start_
      -- CP-element group 190: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Update/cr
      -- 
    cr_3703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(190), ack => type_cast_1491_inst_req_1); -- 
    convTransposeA_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(192) & convTransposeA_CP_3049_elements(212);
      gj_convTransposeA_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	77 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Sample/ra
      -- 
    ra_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1491_inst_ack_0, ack => convTransposeA_CP_3049_elements(191)); -- 
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	210 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1491_Update/ca
      -- 
    ca_3704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1491_inst_ack_1, ack => convTransposeA_CP_3049_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	60 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Sample/rr
      -- 
    rr_3712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(193), ack => type_cast_1515_inst_req_0); -- 
    convTransposeA_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(60) & convTransposeA_CP_3049_elements(195);
      gj_convTransposeA_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: 	200 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_update_start_
      -- CP-element group 194: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Update/cr
      -- 
    cr_3717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(194), ack => type_cast_1515_inst_req_1); -- 
    convTransposeA_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(196) & convTransposeA_CP_3049_elements(200);
      gj_convTransposeA_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	58 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Sample/ra
      -- 
    ra_3713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1515_inst_ack_0, ack => convTransposeA_CP_3049_elements(195)); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	200 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (16) 
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1515_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_resized_1
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_scaled_1
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_computed_1
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_resize_1/$entry
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_resize_1/$exit
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_resize_1/index_resize_req
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_resize_1/index_resize_ack
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_scale_1/$entry
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_scale_1/$exit
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_scale_1/scale_rename_req
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_index_scale_1/scale_rename_ack
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Sample/req
      -- 
    ca_3718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1515_inst_ack_1, ack => convTransposeA_CP_3049_elements(196)); -- 
    req_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(196), ack => array_obj_ref_1521_index_offset_req_0); -- 
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	202 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	202 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_request/req
      -- CP-element group 197: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_request/$entry
      -- 
    req_3758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(197), ack => addr_of_1522_final_reg_req_0); -- 
    convTransposeA_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(201) & convTransposeA_CP_3049_elements(202);
      gj_convTransposeA_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	51 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	203 
    -- CP-element group 198: 	206 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	203 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_complete/$entry
      -- CP-element group 198: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_complete/req
      -- CP-element group 198: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_update_start_
      -- 
    req_3763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(198), ack => addr_of_1522_final_reg_req_1); -- 
    convTransposeA_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(203) & convTransposeA_CP_3049_elements(206);
      gj_convTransposeA_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	51 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	201 
    -- CP-element group 199: 	202 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_update_start
      -- CP-element group 199: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Update/req
      -- 
    req_3748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(199), ack => array_obj_ref_1521_index_offset_req_1); -- 
    convTransposeA_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(201) & convTransposeA_CP_3049_elements(202);
      gj_convTransposeA_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	196 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	277 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	194 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_sample_complete
      -- CP-element group 200: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Sample/ack
      -- 
    ack_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1521_index_offset_ack_0, ack => convTransposeA_CP_3049_elements(200)); -- 
    -- CP-element group 201:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	199 
    -- CP-element group 201:  members (8) 
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_root_address_calculated
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_offset_calculated
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_final_index_sum_regn_Update/ack
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_base_plus_offset/$entry
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_base_plus_offset/$exit
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_base_plus_offset/sum_rename_req
      -- CP-element group 201: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1521_base_plus_offset/sum_rename_ack
      -- 
    ack_3749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1521_index_offset_ack_1, ack => convTransposeA_CP_3049_elements(201)); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	197 
    -- CP-element group 202: successors 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	197 
    -- CP-element group 202: 	199 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_request/ack
      -- CP-element group 202: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_request/$exit
      -- CP-element group 202: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_sample_completed_
      -- 
    ack_3759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1522_final_reg_ack_0, ack => convTransposeA_CP_3049_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	198 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	198 
    -- CP-element group 203:  members (19) 
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_word_addrgen/root_register_req
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_word_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_root_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_address_resized
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_addr_resize/$entry
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_addr_resize/$exit
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_word_addrgen/root_register_ack
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_complete/$exit
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_addr_resize/base_resize_req
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_addr_resize/base_resize_ack
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_plus_offset/$entry
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_complete/ack
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_word_addrgen/$exit
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_word_addrgen/$entry
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_plus_offset/sum_rename_ack
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_plus_offset/sum_rename_req
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_base_plus_offset/$exit
      -- CP-element group 203: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1522_update_completed_
      -- 
    ack_3764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1522_final_reg_ack_1, ack => convTransposeA_CP_3049_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/word_access_start/word_0/rr
      -- CP-element group 204: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/word_access_start/word_0/$entry
      -- CP-element group 204: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/word_access_start/$entry
      -- CP-element group 204: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_sample_start_
      -- 
    rr_3797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(204), ack => ptr_deref_1526_load_0_req_0); -- 
    convTransposeA_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(203) & convTransposeA_CP_3049_elements(206);
      gj_convTransposeA_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: 	222 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_update_start_
      -- CP-element group 205: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/$entry
      -- CP-element group 205: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/word_access_complete/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/word_access_complete/$entry
      -- CP-element group 205: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/word_access_complete/word_0/cr
      -- 
    cr_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(205), ack => ptr_deref_1526_load_0_req_1); -- 
    convTransposeA_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(207) & convTransposeA_CP_3049_elements(222);
      gj_convTransposeA_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	198 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/word_access_start/word_0/ra
      -- CP-element group 206: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_sample_completed_
      -- 
    ra_3798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1526_load_0_ack_0, ack => convTransposeA_CP_3049_elements(206)); -- 
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	220 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/ptr_deref_1526_Merge/merge_ack
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/ptr_deref_1526_Merge/merge_req
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/ptr_deref_1526_Merge/$exit
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/ptr_deref_1526_Merge/$entry
      -- CP-element group 207: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1526_Update/word_access_complete/word_0/ca
      -- 
    ca_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1526_load_0_ack_1, ack => convTransposeA_CP_3049_elements(207)); -- 
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	213 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	214 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	214 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_request/req
      -- CP-element group 208: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_request/$entry
      -- 
    req_3854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(208), ack => addr_of_1545_final_reg_req_0); -- 
    convTransposeA_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(213) & convTransposeA_CP_3049_elements(214);
      gj_convTransposeA_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	51 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	215 
    -- CP-element group 209: 	218 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	215 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_complete/req
      -- CP-element group 209: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_complete/$entry
      -- CP-element group 209: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_update_start_
      -- 
    req_3859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(209), ack => addr_of_1545_final_reg_req_1); -- 
    convTransposeA_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(215) & convTransposeA_CP_3049_elements(218);
      gj_convTransposeA_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	184 
    -- CP-element group 210: 	188 
    -- CP-element group 210: 	192 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (13) 
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Sample/req
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_scale_1/scale_rename_ack
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_scale_1/scale_rename_req
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_scale_1/$exit
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_scale_1/$entry
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_resize_1/index_resize_ack
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_resize_1/index_resize_req
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_resize_1/$exit
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_resize_1/$entry
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_computed_1
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_scaled_1
      -- CP-element group 210: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_index_resized_1
      -- 
    req_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(210), ack => array_obj_ref_1544_index_offset_req_0); -- 
    convTransposeA_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(184) & convTransposeA_CP_3049_elements(188) & convTransposeA_CP_3049_elements(192);
      gj_convTransposeA_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	51 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: 	214 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Update/req
      -- CP-element group 211: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_update_start
      -- 
    req_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(211), ack => array_obj_ref_1544_index_offset_req_1); -- 
    convTransposeA_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(213) & convTransposeA_CP_3049_elements(214);
      gj_convTransposeA_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	277 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	182 
    -- CP-element group 212: 	186 
    -- CP-element group 212: 	190 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Sample/ack
      -- CP-element group 212: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_sample_complete
      -- 
    ack_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1544_index_offset_ack_0, ack => convTransposeA_CP_3049_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	208 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (8) 
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_base_plus_offset/sum_rename_ack
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_base_plus_offset/sum_rename_req
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_base_plus_offset/$exit
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_base_plus_offset/$entry
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Update/ack
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_final_index_sum_regn_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_offset_calculated
      -- CP-element group 213: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/array_obj_ref_1544_root_address_calculated
      -- 
    ack_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1544_index_offset_ack_1, ack => convTransposeA_CP_3049_elements(213)); -- 
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	208 
    -- CP-element group 214: successors 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	208 
    -- CP-element group 214: 	211 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_request/ack
      -- CP-element group 214: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_request/$exit
      -- CP-element group 214: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_sample_completed_
      -- 
    ack_3855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1545_final_reg_ack_0, ack => convTransposeA_CP_3049_elements(214)); -- 
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	209 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	209 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_complete/ack
      -- CP-element group 215: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_complete/$exit
      -- CP-element group 215: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/addr_of_1545_update_completed_
      -- 
    ack_3860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1545_final_reg_ack_1, ack => convTransposeA_CP_3049_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Sample/req
      -- CP-element group 216: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_sample_start_
      -- 
    req_3868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(216), ack => W_arrayidx72_1547_delayed_6_0_1547_inst_req_0); -- 
    convTransposeA_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(215) & convTransposeA_CP_3049_elements(218);
      gj_convTransposeA_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	222 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Update/req
      -- CP-element group 217: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_update_start_
      -- 
    req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(217), ack => W_arrayidx72_1547_delayed_6_0_1547_inst_req_1); -- 
    convTransposeA_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(219) & convTransposeA_CP_3049_elements(222);
      gj_convTransposeA_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	209 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Sample/ack
      -- CP-element group 218: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Sample/$exit
      -- CP-element group 218: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_sample_completed_
      -- 
    ack_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx72_1547_delayed_6_0_1547_inst_ack_0, ack => convTransposeA_CP_3049_elements(218)); -- 
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (19) 
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Update/$exit
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_Update/ack
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_addr_resize/$exit
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_addr_resize/base_resize_req
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_addr_resize/base_resize_ack
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_plus_offset/$entry
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1549_update_completed_
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_addr_resize/$entry
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_address_resized
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_word_addrgen/root_register_ack
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_word_addrgen/root_register_req
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_root_address_calculated
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_word_addrgen/$exit
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_word_addrgen/$entry
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_word_address_calculated
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_plus_offset/sum_rename_ack
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_plus_offset/sum_rename_req
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_address_calculated
      -- CP-element group 219: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_base_plus_offset/$exit
      -- 
    ack_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx72_1547_delayed_6_0_1547_inst_ack_1, ack => convTransposeA_CP_3049_elements(219)); -- 
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	207 
    -- CP-element group 220: 	219 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (9) 
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/word_access_start/word_0/rr
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/word_access_start/word_0/$entry
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/word_access_start/$entry
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/ptr_deref_1551_Split/split_ack
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/ptr_deref_1551_Split/split_req
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/ptr_deref_1551_Split/$exit
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/ptr_deref_1551_Split/$entry
      -- CP-element group 220: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/$entry
      -- 
    rr_3912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(220), ack => ptr_deref_1551_store_0_req_0); -- 
    convTransposeA_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(207) & convTransposeA_CP_3049_elements(219) & convTransposeA_CP_3049_elements(222);
      gj_convTransposeA_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (5) 
      -- CP-element group 221: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_update_start_
      -- CP-element group 221: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/word_access_complete/$entry
      -- CP-element group 221: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/word_access_complete/word_0/$entry
      -- CP-element group 221: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/word_access_complete/word_0/cr
      -- 
    cr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(221), ack => ptr_deref_1551_store_0_req_1); -- 
    convTransposeA_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeA_CP_3049_elements(223);
      gj_convTransposeA_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	205 
    -- CP-element group 222: 	217 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/word_access_start/word_0/ra
      -- CP-element group 222: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_sample_completed_
      -- CP-element group 222: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/word_access_start/word_0/$exit
      -- CP-element group 222: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/word_access_start/$exit
      -- CP-element group 222: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Sample/$exit
      -- 
    ra_3913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1551_store_0_ack_0, ack => convTransposeA_CP_3049_elements(222)); -- 
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	277 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (5) 
      -- CP-element group 223: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/word_access_complete/$exit
      -- CP-element group 223: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/word_access_complete/word_0/$exit
      -- CP-element group 223: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/ptr_deref_1551_Update/word_access_complete/word_0/ca
      -- 
    ca_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1551_store_0_ack_1, ack => convTransposeA_CP_3049_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	123 
    -- CP-element group 224: marked-predecessors 
    -- CP-element group 224: 	226 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_sample_start_
      -- 
    rr_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(224), ack => type_cast_1556_inst_req_0); -- 
    convTransposeA_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(123) & convTransposeA_CP_3049_elements(226);
      gj_convTransposeA_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	54 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: 	242 
    -- CP-element group 225: 	258 
    -- CP-element group 225: 	266 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Update/cr
      -- CP-element group 225: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_update_start_
      -- 
    cr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(225), ack => type_cast_1556_inst_req_1); -- 
    convTransposeA_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(227) & convTransposeA_CP_3049_elements(242) & convTransposeA_CP_3049_elements(258) & convTransposeA_CP_3049_elements(266);
      gj_convTransposeA_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	119 
    -- CP-element group 226: 	224 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Sample/ra
      -- CP-element group 226: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_sample_completed_
      -- 
    ra_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1556_inst_ack_0, ack => convTransposeA_CP_3049_elements(226)); -- 
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	240 
    -- CP-element group 227: 	256 
    -- CP-element group 227: 	264 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	118 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Update/ca
      -- CP-element group 227: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1556_update_completed_
      -- 
    ca_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1556_inst_ack_1, ack => convTransposeA_CP_3049_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	51 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_sample_start_
      -- 
    rr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(228), ack => type_cast_1560_inst_req_0); -- 
    convTransposeA_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(51) & convTransposeA_CP_3049_elements(230);
      gj_convTransposeA_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	54 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: 	242 
    -- CP-element group 229: 	258 
    -- CP-element group 229: 	266 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_update_start_
      -- 
    cr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(229), ack => type_cast_1560_inst_req_1); -- 
    convTransposeA_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(231) & convTransposeA_CP_3049_elements(242) & convTransposeA_CP_3049_elements(258) & convTransposeA_CP_3049_elements(266);
      gj_convTransposeA_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Sample/ra
      -- CP-element group 230: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_sample_completed_
      -- 
    ra_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1560_inst_ack_0, ack => convTransposeA_CP_3049_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	240 
    -- CP-element group 231: 	256 
    -- CP-element group 231: 	264 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	118 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Update/ca
      -- CP-element group 231: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1560_update_completed_
      -- 
    ca_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1560_inst_ack_1, ack => convTransposeA_CP_3049_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	102 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	234 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_sample_start_
      -- 
    req_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(232), ack => W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_req_0); -- 
    convTransposeA_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(102) & convTransposeA_CP_3049_elements(234);
      gj_convTransposeA_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: 	258 
    -- CP-element group 233: 	266 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_update_start_
      -- CP-element group 233: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Update/req
      -- 
    req_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(233), ack => W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_req_1); -- 
    convTransposeA_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(235) & convTransposeA_CP_3049_elements(258) & convTransposeA_CP_3049_elements(266);
      gj_convTransposeA_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	98 
    -- CP-element group 234: 	232 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Sample/ack
      -- CP-element group 234: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_sample_completed_
      -- 
    ack_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_ack_0, ack => convTransposeA_CP_3049_elements(234)); -- 
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	256 
    -- CP-element group 235: 	264 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1583_Update/ack
      -- 
    ack_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_ack_1, ack => convTransposeA_CP_3049_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	123 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_sample_start_
      -- 
    req_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(236), ack => W_add87_1582_delayed_1_0_1589_inst_req_0); -- 
    convTransposeA_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(123) & convTransposeA_CP_3049_elements(238);
      gj_convTransposeA_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	54 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Update/req
      -- CP-element group 237: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_update_start_
      -- 
    req_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(237), ack => W_add87_1582_delayed_1_0_1589_inst_req_1); -- 
    convTransposeA_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(239);
      gj_convTransposeA_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	119 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Sample/ack
      -- CP-element group 238: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_sample_completed_
      -- 
    ack_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add87_1582_delayed_1_0_1589_inst_ack_0, ack => convTransposeA_CP_3049_elements(238)); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	277 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	118 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Update/ack
      -- CP-element group 239: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1591_update_completed_
      -- 
    ack_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add87_1582_delayed_1_0_1589_inst_ack_1, ack => convTransposeA_CP_3049_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	227 
    -- CP-element group 240: 	231 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Sample/rr
      -- CP-element group 240: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_sample_start_
      -- 
    rr_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(240), ack => type_cast_1601_inst_req_0); -- 
    convTransposeA_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(227) & convTransposeA_CP_3049_elements(231) & convTransposeA_CP_3049_elements(242);
      gj_convTransposeA_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	54 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: 	274 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_update_start_
      -- CP-element group 241: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Update/cr
      -- CP-element group 241: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Update/$entry
      -- 
    cr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(241), ack => type_cast_1601_inst_req_1); -- 
    convTransposeA_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(243) & convTransposeA_CP_3049_elements(274);
      gj_convTransposeA_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	225 
    -- CP-element group 242: 	229 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Sample/ra
      -- 
    ra_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_0, ack => convTransposeA_CP_3049_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	272 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	76 
    -- CP-element group 243: 	97 
    -- CP-element group 243: 	139 
    -- CP-element group 243: 	160 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Update/ca
      -- CP-element group 243: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1601_Update/$exit
      -- 
    ca_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_1, ack => convTransposeA_CP_3049_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	144 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_sample_start_
      -- 
    req_4002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(244), ack => W_input_dim1x_x1_1599_delayed_2_0_1609_inst_req_0); -- 
    convTransposeA_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(144) & convTransposeA_CP_3049_elements(246);
      gj_convTransposeA_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	54 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	274 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Update/req
      -- CP-element group 245: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_update_start_
      -- 
    req_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(245), ack => W_input_dim1x_x1_1599_delayed_2_0_1609_inst_req_1); -- 
    convTransposeA_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(247) & convTransposeA_CP_3049_elements(274);
      gj_convTransposeA_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	140 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Sample/ack
      -- CP-element group 246: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_sample_completed_
      -- 
    ack_4003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_1599_delayed_2_0_1609_inst_ack_0, ack => convTransposeA_CP_3049_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	272 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	76 
    -- CP-element group 247: 	97 
    -- CP-element group 247: 	139 
    -- CP-element group 247: 	160 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Update/ack
      -- CP-element group 247: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1611_update_completed_
      -- 
    ack_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_1599_delayed_2_0_1609_inst_ack_1, ack => convTransposeA_CP_3049_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	165 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Sample/$entry
      -- 
    req_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(248), ack => W_input_dim0x_x1_1619_delayed_2_0_1632_inst_req_0); -- 
    convTransposeA_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(165) & convTransposeA_CP_3049_elements(250);
      gj_convTransposeA_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	54 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	274 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Update/req
      -- CP-element group 249: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_update_start_
      -- 
    req_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(249), ack => W_input_dim0x_x1_1619_delayed_2_0_1632_inst_req_1); -- 
    convTransposeA_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(251) & convTransposeA_CP_3049_elements(274);
      gj_convTransposeA_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	161 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Sample/ack
      -- CP-element group 250: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Sample/$exit
      -- 
    ack_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_1619_delayed_2_0_1632_inst_ack_0, ack => convTransposeA_CP_3049_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	272 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	160 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Update/ack
      -- CP-element group 251: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1634_update_completed_
      -- 
    ack_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_1619_delayed_2_0_1632_inst_ack_1, ack => convTransposeA_CP_3049_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	81 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_sample_start_
      -- 
    req_4030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(252), ack => W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_req_0); -- 
    convTransposeA_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(81) & convTransposeA_CP_3049_elements(254);
      gj_convTransposeA_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	54 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Update/req
      -- CP-element group 253: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_update_start_
      -- 
    req_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(253), ack => W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_req_1); -- 
    convTransposeA_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(255);
      gj_convTransposeA_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	77 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Sample/ack
      -- CP-element group 254: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_sample_completed_
      -- 
    ack_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_ack_0, ack => convTransposeA_CP_3049_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	277 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	76 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Update/ack
      -- CP-element group 255: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1644_update_completed_
      -- 
    ack_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_ack_1, ack => convTransposeA_CP_3049_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	227 
    -- CP-element group 256: 	231 
    -- CP-element group 256: 	235 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_sample_start_
      -- 
    req_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(256), ack => W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_req_0); -- 
    convTransposeA_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(227) & convTransposeA_CP_3049_elements(231) & convTransposeA_CP_3049_elements(235) & convTransposeA_CP_3049_elements(258);
      gj_convTransposeA_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	54 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Update/req
      -- CP-element group 257: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_update_start_
      -- 
    req_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(257), ack => W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_req_1); -- 
    convTransposeA_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(259);
      gj_convTransposeA_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	225 
    -- CP-element group 258: 	229 
    -- CP-element group 258: 	233 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Sample/ack
      -- CP-element group 258: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_sample_completed_
      -- 
    ack_4045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_ack_0, ack => convTransposeA_CP_3049_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	277 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	97 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Update/ack
      -- CP-element group 259: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/assign_stmt_1653_update_completed_
      -- 
    ack_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_ack_1, ack => convTransposeA_CP_3049_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	81 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_sample_start_
      -- 
    rr_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(260), ack => type_cast_1665_inst_req_0); -- 
    convTransposeA_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(81) & convTransposeA_CP_3049_elements(262);
      gj_convTransposeA_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	54 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_update_start_
      -- 
    cr_4063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(261), ack => type_cast_1665_inst_req_1); -- 
    convTransposeA_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(263);
      gj_convTransposeA_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	77 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Sample/ra
      -- CP-element group 262: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_sample_completed_
      -- 
    ra_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_0, ack => convTransposeA_CP_3049_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	277 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	76 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1665_update_completed_
      -- 
    ca_4064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_1, ack => convTransposeA_CP_3049_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	227 
    -- CP-element group 264: 	231 
    -- CP-element group 264: 	235 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Sample/rr
      -- CP-element group 264: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Sample/$entry
      -- 
    rr_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(264), ack => type_cast_1680_inst_req_0); -- 
    convTransposeA_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(227) & convTransposeA_CP_3049_elements(231) & convTransposeA_CP_3049_elements(235) & convTransposeA_CP_3049_elements(266);
      gj_convTransposeA_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	54 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_update_start_
      -- CP-element group 265: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Update/cr
      -- CP-element group 265: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Update/$entry
      -- 
    cr_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(265), ack => type_cast_1680_inst_req_1); -- 
    convTransposeA_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(267);
      gj_convTransposeA_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	225 
    -- CP-element group 266: 	229 
    -- CP-element group 266: 	233 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Sample/ra
      -- 
    ra_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1680_inst_ack_0, ack => convTransposeA_CP_3049_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	277 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	97 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Update/ca
      -- CP-element group 267: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1680_Update/$exit
      -- 
    ca_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1680_inst_ack_1, ack => convTransposeA_CP_3049_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	165 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Sample/$entry
      -- 
    rr_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(268), ack => type_cast_1708_inst_req_0); -- 
    convTransposeA_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(165) & convTransposeA_CP_3049_elements(270);
      gj_convTransposeA_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	54 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	274 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Update/cr
      -- CP-element group 269: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_update_start_
      -- 
    cr_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(269), ack => type_cast_1708_inst_req_1); -- 
    convTransposeA_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(271) & convTransposeA_CP_3049_elements(274);
      gj_convTransposeA_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	161 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Sample/ra
      -- CP-element group 270: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Sample/$exit
      -- 
    ra_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1708_inst_ack_0, ack => convTransposeA_CP_3049_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	160 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_Update/ca
      -- CP-element group 271: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1708_update_completed_
      -- 
    ca_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1708_inst_ack_1, ack => convTransposeA_CP_3049_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	243 
    -- CP-element group 272: 	247 
    -- CP-element group 272: 	251 
    -- CP-element group 272: 	271 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Sample/rr
      -- 
    rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(272), ack => type_cast_1723_inst_req_0); -- 
    convTransposeA_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(243) & convTransposeA_CP_3049_elements(247) & convTransposeA_CP_3049_elements(251) & convTransposeA_CP_3049_elements(271) & convTransposeA_CP_3049_elements(274);
      gj_convTransposeA_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_update_start_
      -- 
    cr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(273), ack => type_cast_1723_inst_req_1); -- 
    convTransposeA_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeA_CP_3049_elements(275);
      gj_convTransposeA_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	241 
    -- CP-element group 274: 	245 
    -- CP-element group 274: 	249 
    -- CP-element group 274: 	269 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Sample/ra
      -- CP-element group 274: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Sample/$exit
      -- 
    ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_0, ack => convTransposeA_CP_3049_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	52 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/type_cast_1723_Update/$exit
      -- 
    ca_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_1, ack => convTransposeA_CP_3049_elements(275)); -- 
    -- CP-element group 276:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	51 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	52 
    -- CP-element group 276:  members (1) 
      -- CP-element group 276: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convTransposeA_CP_3049_elements(276) is a control-delay.
    cp_element_276_delay: control_delay_element  generic map(name => " 276_delay", delay_value => 1)  port map(req => convTransposeA_CP_3049_elements(51), ack => convTransposeA_CP_3049_elements(276), clk => clk, reset =>reset);
    -- CP-element group 277:  join  transition  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	54 
    -- CP-element group 277: 	200 
    -- CP-element group 277: 	212 
    -- CP-element group 277: 	223 
    -- CP-element group 277: 	239 
    -- CP-element group 277: 	255 
    -- CP-element group 277: 	259 
    -- CP-element group 277: 	263 
    -- CP-element group 277: 	267 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	48 
    -- CP-element group 277:  members (1) 
      -- CP-element group 277: 	 branch_block_stmt_1298/do_while_stmt_1443/do_while_stmt_1443_loop_body/$exit
      -- 
    convTransposeA_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(54) & convTransposeA_CP_3049_elements(200) & convTransposeA_CP_3049_elements(212) & convTransposeA_CP_3049_elements(223) & convTransposeA_CP_3049_elements(239) & convTransposeA_CP_3049_elements(255) & convTransposeA_CP_3049_elements(259) & convTransposeA_CP_3049_elements(263) & convTransposeA_CP_3049_elements(267);
      gj_convTransposeA_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	47 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_exit/$exit
      -- CP-element group 278: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_exit/ack
      -- 
    ack_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1443_branch_ack_0, ack => convTransposeA_CP_3049_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	47 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (2) 
      -- CP-element group 279: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_taken/ack
      -- CP-element group 279: 	 branch_block_stmt_1298/do_while_stmt_1443/loop_taken/$exit
      -- 
    ack_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1443_branch_ack_1, ack => convTransposeA_CP_3049_elements(279)); -- 
    -- CP-element group 280:  transition  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	45 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	1 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_1298/do_while_stmt_1443/$exit
      -- 
    convTransposeA_CP_3049_elements(280) <= convTransposeA_CP_3049_elements(45);
    -- CP-element group 281:  merge  transition  place  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	1 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (15) 
      -- CP-element group 281: 	 branch_block_stmt_1298/merge_stmt_1746__exit__
      -- CP-element group 281: 	 branch_block_stmt_1298/assign_stmt_1751__entry__
      -- CP-element group 281: 	 branch_block_stmt_1298/if_stmt_1742_if_link/$exit
      -- CP-element group 281: 	 branch_block_stmt_1298/if_stmt_1742_if_link/if_choice_transition
      -- CP-element group 281: 	 branch_block_stmt_1298/ifx_xend122_whilex_xend
      -- CP-element group 281: 	 branch_block_stmt_1298/assign_stmt_1751/$entry
      -- CP-element group 281: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Sample/req
      -- CP-element group 281: 	 branch_block_stmt_1298/ifx_xend122_whilex_xend_PhiReq/$entry
      -- CP-element group 281: 	 branch_block_stmt_1298/ifx_xend122_whilex_xend_PhiReq/$exit
      -- CP-element group 281: 	 branch_block_stmt_1298/merge_stmt_1746_PhiReqMerge
      -- CP-element group 281: 	 branch_block_stmt_1298/merge_stmt_1746_PhiAck/$entry
      -- CP-element group 281: 	 branch_block_stmt_1298/merge_stmt_1746_PhiAck/$exit
      -- CP-element group 281: 	 branch_block_stmt_1298/merge_stmt_1746_PhiAck/dummy
      -- 
    if_choice_transition_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1742_branch_ack_1, ack => convTransposeA_CP_3049_elements(281)); -- 
    req_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(281), ack => WPIPE_Block0_done_1748_inst_req_0); -- 
    -- CP-element group 282:  merge  transition  place  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	1 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (5) 
      -- CP-element group 282: 	 branch_block_stmt_1298/if_stmt_1742__exit__
      -- CP-element group 282: 	 branch_block_stmt_1298/merge_stmt_1746__entry__
      -- CP-element group 282: 	 branch_block_stmt_1298/if_stmt_1742_else_link/$exit
      -- CP-element group 282: 	 branch_block_stmt_1298/if_stmt_1742_else_link/else_choice_transition
      -- CP-element group 282: 	 branch_block_stmt_1298/merge_stmt_1746_dead_link/$entry
      -- 
    else_choice_transition_4133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1742_branch_ack_0, ack => convTransposeA_CP_3049_elements(282)); -- 
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Sample/ack
      -- CP-element group 283: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Update/req
      -- 
    ack_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1748_inst_ack_0, ack => convTransposeA_CP_3049_elements(283)); -- 
    req_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(283), ack => WPIPE_Block0_done_1748_inst_req_1); -- 
    -- CP-element group 284:  transition  place  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (16) 
      -- CP-element group 284: 	 $exit
      -- CP-element group 284: 	 branch_block_stmt_1298/$exit
      -- CP-element group 284: 	 branch_block_stmt_1298/branch_block_stmt_1298__exit__
      -- CP-element group 284: 	 branch_block_stmt_1298/assign_stmt_1751__exit__
      -- CP-element group 284: 	 branch_block_stmt_1298/return__
      -- CP-element group 284: 	 branch_block_stmt_1298/merge_stmt_1753__exit__
      -- CP-element group 284: 	 branch_block_stmt_1298/assign_stmt_1751/$exit
      -- CP-element group 284: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_1298/assign_stmt_1751/WPIPE_Block0_done_1748_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_1298/return___PhiReq/$entry
      -- CP-element group 284: 	 branch_block_stmt_1298/return___PhiReq/$exit
      -- CP-element group 284: 	 branch_block_stmt_1298/merge_stmt_1753_PhiReqMerge
      -- CP-element group 284: 	 branch_block_stmt_1298/merge_stmt_1753_PhiAck/$entry
      -- CP-element group 284: 	 branch_block_stmt_1298/merge_stmt_1753_PhiAck/$exit
      -- CP-element group 284: 	 branch_block_stmt_1298/merge_stmt_1753_PhiAck/dummy
      -- 
    ack_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1748_inst_ack_1, ack => convTransposeA_CP_3049_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	43 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Sample/ra
      -- 
    ra_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_0, ack => convTransposeA_CP_3049_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	43 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/Update/ca
      -- 
    ca_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_1, ack => convTransposeA_CP_3049_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	291 
    -- CP-element group 287:  members (5) 
      -- CP-element group 287: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 287: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 287: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/$exit
      -- CP-element group 287: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1426/SplitProtocol/$exit
      -- CP-element group 287: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_4177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_4177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(287), ack => phi_stmt_1423_req_0); -- 
    convTransposeA_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(285) & convTransposeA_CP_3049_elements(286);
      gj_convTransposeA_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	43 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Sample/ra
      -- 
    ra_4194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_0, ack => convTransposeA_CP_3049_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	43 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/Update/ca
      -- 
    ca_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_1, ack => convTransposeA_CP_3049_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (5) 
      -- CP-element group 290: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/$exit
      -- CP-element group 290: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/$exit
      -- CP-element group 290: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1422/SplitProtocol/$exit
      -- CP-element group 290: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/phi_stmt_1419/phi_stmt_1419_req
      -- 
    phi_stmt_1419_req_4200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1419_req_4200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3049_elements(290), ack => phi_stmt_1419_req_0); -- 
    convTransposeA_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(288) & convTransposeA_CP_3049_elements(289);
      gj_convTransposeA_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  fork  transition  place  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	287 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_1298/entry_whilex_xbody_PhiReq/$exit
      -- CP-element group 291: 	 branch_block_stmt_1298/merge_stmt_1413_PhiReqMerge
      -- CP-element group 291: 	 branch_block_stmt_1298/merge_stmt_1413_PhiAck/$entry
      -- 
    convTransposeA_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(287) & convTransposeA_CP_3049_elements(290);
      gj_convTransposeA_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (1) 
      -- CP-element group 292: 	 branch_block_stmt_1298/merge_stmt_1413_PhiAck/phi_stmt_1419_ack
      -- 
    phi_stmt_1419_ack_4205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1419_ack_0, ack => convTransposeA_CP_3049_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (1) 
      -- CP-element group 293: 	 branch_block_stmt_1298/merge_stmt_1413_PhiAck/phi_stmt_1423_ack
      -- 
    phi_stmt_1423_ack_4206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1423_ack_0, ack => convTransposeA_CP_3049_elements(293)); -- 
    -- CP-element group 294:  join  transition  place  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	44 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_1298/merge_stmt_1413__exit__
      -- CP-element group 294: 	 branch_block_stmt_1298/do_while_stmt_1443__entry__
      -- CP-element group 294: 	 branch_block_stmt_1298/merge_stmt_1413_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3049_elements(292) & convTransposeA_CP_3049_elements(293);
      gj_convTransposeA_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3049_elements(294), clk => clk, reset => reset); --
    end block;
    convTransposeA_do_while_stmt_1443_terminator_4116: loop_terminator -- 
      generic map (name => " convTransposeA_do_while_stmt_1443_terminator_4116", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convTransposeA_CP_3049_elements(48),loop_continue => convTransposeA_CP_3049_elements(279),loop_terminate => convTransposeA_CP_3049_elements(278),loop_back => convTransposeA_CP_3049_elements(46),loop_exit => convTransposeA_CP_3049_elements(45),clk => clk, reset => reset); -- 
    phi_stmt_1445_phi_seq_3422_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3049_elements(63);
      convTransposeA_CP_3049_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3049_elements(66);
      convTransposeA_CP_3049_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3049_elements(68);
      convTransposeA_CP_3049_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3049_elements(61);
      convTransposeA_CP_3049_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3049_elements(74);
      convTransposeA_CP_3049_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3049_elements(75);
      convTransposeA_CP_3049_elements(62) <= phi_mux_reqs(1);
      phi_stmt_1445_phi_seq_3422 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1445_phi_seq_3422") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3049_elements(53), 
          phi_sample_ack => convTransposeA_CP_3049_elements(59), 
          phi_update_req => convTransposeA_CP_3049_elements(55), 
          phi_update_ack => convTransposeA_CP_3049_elements(60), 
          phi_mux_ack => convTransposeA_CP_3049_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1450_phi_seq_3476_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3049_elements(82);
      convTransposeA_CP_3049_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3049_elements(91);
      convTransposeA_CP_3049_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3049_elements(92);
      convTransposeA_CP_3049_elements(83) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3049_elements(84);
      convTransposeA_CP_3049_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3049_elements(95);
      convTransposeA_CP_3049_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3049_elements(96);
      convTransposeA_CP_3049_elements(85) <= phi_mux_reqs(1);
      phi_stmt_1450_phi_seq_3476 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1450_phi_seq_3476") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3049_elements(78), 
          phi_sample_ack => convTransposeA_CP_3049_elements(79), 
          phi_update_req => convTransposeA_CP_3049_elements(80), 
          phi_update_ack => convTransposeA_CP_3049_elements(81), 
          phi_mux_ack => convTransposeA_CP_3049_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1455_phi_seq_3530_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3049_elements(103);
      convTransposeA_CP_3049_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3049_elements(112);
      convTransposeA_CP_3049_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3049_elements(113);
      convTransposeA_CP_3049_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3049_elements(105);
      convTransposeA_CP_3049_elements(114)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3049_elements(116);
      convTransposeA_CP_3049_elements(115)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3049_elements(117);
      convTransposeA_CP_3049_elements(106) <= phi_mux_reqs(1);
      phi_stmt_1455_phi_seq_3530 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1455_phi_seq_3530") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3049_elements(99), 
          phi_sample_ack => convTransposeA_CP_3049_elements(100), 
          phi_update_req => convTransposeA_CP_3049_elements(101), 
          phi_update_ack => convTransposeA_CP_3049_elements(102), 
          phi_mux_ack => convTransposeA_CP_3049_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1460_phi_seq_3574_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3049_elements(124);
      convTransposeA_CP_3049_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3049_elements(133);
      convTransposeA_CP_3049_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3049_elements(134);
      convTransposeA_CP_3049_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3049_elements(126);
      convTransposeA_CP_3049_elements(135)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3049_elements(135);
      convTransposeA_CP_3049_elements(136)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3049_elements(137);
      convTransposeA_CP_3049_elements(127) <= phi_mux_reqs(1);
      phi_stmt_1460_phi_seq_3574 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1460_phi_seq_3574") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3049_elements(120), 
          phi_sample_ack => convTransposeA_CP_3049_elements(121), 
          phi_update_req => convTransposeA_CP_3049_elements(122), 
          phi_update_ack => convTransposeA_CP_3049_elements(123), 
          phi_mux_ack => convTransposeA_CP_3049_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1465_phi_seq_3618_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3049_elements(145);
      convTransposeA_CP_3049_elements(150)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3049_elements(154);
      convTransposeA_CP_3049_elements(151)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3049_elements(155);
      convTransposeA_CP_3049_elements(146) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3049_elements(147);
      convTransposeA_CP_3049_elements(156)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3049_elements(156);
      convTransposeA_CP_3049_elements(157)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3049_elements(158);
      convTransposeA_CP_3049_elements(148) <= phi_mux_reqs(1);
      phi_stmt_1465_phi_seq_3618 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1465_phi_seq_3618") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3049_elements(141), 
          phi_sample_ack => convTransposeA_CP_3049_elements(142), 
          phi_update_req => convTransposeA_CP_3049_elements(143), 
          phi_update_ack => convTransposeA_CP_3049_elements(144), 
          phi_mux_ack => convTransposeA_CP_3049_elements(149), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1470_phi_seq_3662_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3049_elements(166);
      convTransposeA_CP_3049_elements(171)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3049_elements(175);
      convTransposeA_CP_3049_elements(172)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3049_elements(176);
      convTransposeA_CP_3049_elements(167) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3049_elements(168);
      convTransposeA_CP_3049_elements(177)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3049_elements(177);
      convTransposeA_CP_3049_elements(178)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3049_elements(179);
      convTransposeA_CP_3049_elements(169) <= phi_mux_reqs(1);
      phi_stmt_1470_phi_seq_3662 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1470_phi_seq_3662") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3049_elements(162), 
          phi_sample_ack => convTransposeA_CP_3049_elements(163), 
          phi_update_req => convTransposeA_CP_3049_elements(164), 
          phi_update_ack => convTransposeA_CP_3049_elements(165), 
          phi_mux_ack => convTransposeA_CP_3049_elements(170), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3374_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convTransposeA_CP_3049_elements(49);
        preds(1)  <= convTransposeA_CP_3049_elements(50);
        entry_tmerge_3374 : transition_merge -- 
          generic map(name => " entry_tmerge_3374")
          port map (preds => preds, symbol_out => convTransposeA_CP_3049_elements(51));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_1675_wire : std_logic_vector(15 downto 0);
    signal MUX_1690_wire : std_logic_vector(15 downto 0);
    signal MUX_1703_wire : std_logic_vector(15 downto 0);
    signal MUX_1718_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1741_wire : std_logic_vector(0 downto 0);
    signal R_idxprom71_1543_resized : std_logic_vector(13 downto 0);
    signal R_idxprom71_1543_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1520_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1520_scaled : std_logic_vector(13 downto 0);
    signal add110_1650 : std_logic_vector(15 downto 0);
    signal add30_1366 : std_logic_vector(15 downto 0);
    signal add64_1502 : std_logic_vector(63 downto 0);
    signal add66_1512 : std_logic_vector(63 downto 0);
    signal add87_1573 : std_logic_vector(15 downto 0);
    signal add87_1582_delayed_1_0_1591 : std_logic_vector(15 downto 0);
    signal add94_1580 : std_logic_vector(15 downto 0);
    signal add_1350 : std_logic_vector(31 downto 0);
    signal add_dest_dim0x_x0_1677 : std_logic_vector(15 downto 0);
    signal add_dest_dim0x_x1_1450 : std_logic_vector(15 downto 0);
    signal add_dest_dim0x_x1_1626_delayed_2_0_1644 : std_logic_vector(15 downto 0);
    signal add_dest_dim0x_x1_at_entry_1419 : std_logic_vector(15 downto 0);
    signal add_dest_dim0x_x1_at_entry_1419_1454_buffered : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x0_1588 : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x0_1632_delayed_1_0_1653 : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x1_1455 : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x1_1577_delayed_1_0_1583 : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x1_at_entry_1423 : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x1_at_entry_1423_1459_buffered : std_logic_vector(15 downto 0);
    signal add_dest_dim1x_x2_1692 : std_logic_vector(15 downto 0);
    signal add_src_0x_x0_1480 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1521_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1521_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1521_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1521_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1521_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1521_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1544_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1544_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1544_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1544_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1544_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1544_root_address : std_logic_vector(13 downto 0);
    signal arrayidx68_1523 : std_logic_vector(31 downto 0);
    signal arrayidx72_1546 : std_logic_vector(31 downto 0);
    signal arrayidx72_1547_delayed_6_0_1549 : std_logic_vector(31 downto 0);
    signal call11_1319 : std_logic_vector(15 downto 0);
    signal call13_1322 : std_logic_vector(15 downto 0);
    signal call14_1325 : std_logic_vector(15 downto 0);
    signal call15_1328 : std_logic_vector(15 downto 0);
    signal call16_1341 : std_logic_vector(15 downto 0);
    signal call18_1353 : std_logic_vector(15 downto 0);
    signal call1_1304 : std_logic_vector(15 downto 0);
    signal call20_1356 : std_logic_vector(15 downto 0);
    signal call22_1359 : std_logic_vector(15 downto 0);
    signal call3_1307 : std_logic_vector(15 downto 0);
    signal call5_1310 : std_logic_vector(15 downto 0);
    signal call7_1313 : std_logic_vector(15 downto 0);
    signal call9_1316 : std_logic_vector(15 downto 0);
    signal call_1301 : std_logic_vector(15 downto 0);
    signal cmp101_1621 : std_logic_vector(0 downto 0);
    signal cmp129_1729 : std_logic_vector(0 downto 0);
    signal cmp_1567 : std_logic_vector(0 downto 0);
    signal conv124_1724 : std_logic_vector(31 downto 0);
    signal conv127_1405 : std_logic_vector(31 downto 0);
    signal conv17_1345 : std_logic_vector(31 downto 0);
    signal conv53_1484 : std_logic_vector(63 downto 0);
    signal conv56_1380 : std_logic_vector(63 downto 0);
    signal conv58_1488 : std_logic_vector(63 downto 0);
    signal conv61_1384 : std_logic_vector(63 downto 0);
    signal conv63_1492 : std_logic_vector(63 downto 0);
    signal conv81_1557 : std_logic_vector(31 downto 0);
    signal conv83_1396 : std_logic_vector(31 downto 0);
    signal conv_1332 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1602 : std_logic_vector(15 downto 0);
    signal idxprom71_1539 : std_logic_vector(63 downto 0);
    signal idxprom_1516 : std_logic_vector(63 downto 0);
    signal ifx_xend122_whilex_xend_taken_1738 : std_logic_vector(0 downto 0);
    signal ifx_xthen103_exec_guard_1631 : std_logic_vector(0 downto 0);
    signal ifx_xthen103_ifx_xend122_taken_1662 : std_logic_vector(0 downto 0);
    signal inc105_1641 : std_logic_vector(15 downto 0);
    signal inc_1608 : std_logic_vector(15 downto 0);
    signal indvar_1445 : std_logic_vector(31 downto 0);
    signal indvar_at_entry_1414 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1735 : std_logic_vector(31 downto 0);
    signal input_dim0x_x0_1720 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_1470 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_1619_delayed_2_0_1634 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_1437 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0_1616 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1465 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1599_delayed_2_0_1611 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_at_entry_1432 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1705 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0_1598 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1460 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_at_entry_1427 : std_logic_vector(15 downto 0);
    signal mul117_1401 : std_logic_vector(15 downto 0);
    signal mul65_1507 : std_logic_vector(63 downto 0);
    signal mul_1497 : std_logic_vector(63 downto 0);
    signal ptr_deref_1526_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1526_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1526_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1526_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1526_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1551_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1551_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1338 : std_logic_vector(31 downto 0);
    signal shr128142_1411 : std_logic_vector(31 downto 0);
    signal shr_1533 : std_logic_vector(63 downto 0);
    signal sub120_1659 : std_logic_vector(15 downto 0);
    signal sub45_1376 : std_logic_vector(15 downto 0);
    signal sub77_1390 : std_logic_vector(15 downto 0);
    signal sub_1371 : std_logic_vector(15 downto 0);
    signal tmp69_1527 : std_logic_vector(63 downto 0);
    signal type_cast_1336_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1364_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1394_wire : std_logic_vector(31 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1422_wire : std_logic_vector(15 downto 0);
    signal type_cast_1426_wire : std_logic_vector(15 downto 0);
    signal type_cast_1449_wire : std_logic_vector(31 downto 0);
    signal type_cast_1453_wire : std_logic_vector(15 downto 0);
    signal type_cast_1458_wire : std_logic_vector(15 downto 0);
    signal type_cast_1463_wire : std_logic_vector(15 downto 0);
    signal type_cast_1468_wire : std_logic_vector(15 downto 0);
    signal type_cast_1473_wire : std_logic_vector(15 downto 0);
    signal type_cast_1531_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1537_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1559_1559_delayed_2_0_1561 : std_logic_vector(31 downto 0);
    signal type_cast_1564_wire : std_logic_vector(31 downto 0);
    signal type_cast_1571_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1577_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1596_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1606_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1639_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1645_1645_delayed_2_0_1666 : std_logic_vector(15 downto 0);
    signal type_cast_1657_1657_delayed_1_0_1681 : std_logic_vector(15 downto 0);
    signal type_cast_1670_wire : std_logic_vector(15 downto 0);
    signal type_cast_1674_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1682_1682_delayed_2_0_1709 : std_logic_vector(15 downto 0);
    signal type_cast_1685_wire : std_logic_vector(15 downto 0);
    signal type_cast_1689_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1697_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1700_wire : std_logic_vector(15 downto 0);
    signal type_cast_1702_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1713_wire : std_logic_vector(15 downto 0);
    signal type_cast_1717_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1733_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1750_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_ifx_xend122_taken_1628 : std_logic_vector(0 downto 0);
    signal whilex_xbody_ifx_xthen103_taken_1624 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_1521_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1521_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1521_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1521_resized_base_address <= "00000000000000";
    array_obj_ref_1544_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1544_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1544_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1544_resized_base_address <= "00000000000000";
    indvar_at_entry_1414 <= "00000000000000000000000000000000";
    input_dim0x_x1_at_entry_1437 <= "0000000000000000";
    input_dim1x_x1_at_entry_1432 <= "0000000000000000";
    input_dim2x_x1_at_entry_1427 <= "0000000000000000";
    ptr_deref_1526_word_offset_0 <= "00000000000000";
    ptr_deref_1551_word_offset_0 <= "00000000000000";
    type_cast_1336_wire_constant <= "00000000000000000000000000010000";
    type_cast_1364_wire_constant <= "0000000000000001";
    type_cast_1388_wire_constant <= "1111111111111100";
    type_cast_1409_wire_constant <= "00000000000000000000000000000010";
    type_cast_1531_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1537_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1571_wire_constant <= "0000000000000100";
    type_cast_1577_wire_constant <= "0000000000000000";
    type_cast_1596_wire_constant <= "0000000000000000";
    type_cast_1606_wire_constant <= "0000000000000001";
    type_cast_1639_wire_constant <= "0000000000000001";
    type_cast_1674_wire_constant <= "0000000000000000";
    type_cast_1689_wire_constant <= "0000000000000000";
    type_cast_1697_wire_constant <= "0000000000000000";
    type_cast_1702_wire_constant <= "0000000000000000";
    type_cast_1717_wire_constant <= "0000000000000000";
    type_cast_1733_wire_constant <= "00000000000000000000000000000001";
    type_cast_1750_wire_constant <= "0000000000000001";
    phi_stmt_1419: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1422_wire;
      req(0) <= phi_stmt_1419_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1419",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1419_ack_0,
          idata => idata,
          odata => add_dest_dim0x_x1_at_entry_1419,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1419
    phi_stmt_1423: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1426_wire;
      req(0) <= phi_stmt_1423_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1423",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1423_ack_0,
          idata => idata,
          odata => add_dest_dim1x_x1_at_entry_1423,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1423
    phi_stmt_1445: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= indvar_at_entry_1414 & type_cast_1449_wire;
      req <= phi_stmt_1445_req_0 & phi_stmt_1445_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1445",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1445_ack_0,
          idata => idata,
          odata => indvar_1445,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1445
    phi_stmt_1450: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1453_wire & add_dest_dim0x_x1_at_entry_1419_1454_buffered;
      req <= phi_stmt_1450_req_0 & phi_stmt_1450_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1450",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1450_ack_0,
          idata => idata,
          odata => add_dest_dim0x_x1_1450,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1450
    phi_stmt_1455: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1458_wire & add_dest_dim1x_x1_at_entry_1423_1459_buffered;
      req <= phi_stmt_1455_req_0 & phi_stmt_1455_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1455",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1455_ack_0,
          idata => idata,
          odata => add_dest_dim1x_x1_1455,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1455
    phi_stmt_1460: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1463_wire & input_dim2x_x1_at_entry_1427;
      req <= phi_stmt_1460_req_0 & phi_stmt_1460_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1460",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1460_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1460,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1460
    phi_stmt_1465: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1468_wire & input_dim1x_x1_at_entry_1432;
      req <= phi_stmt_1465_req_0 & phi_stmt_1465_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1465",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1465_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1465,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1465
    phi_stmt_1470: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1473_wire & input_dim0x_x1_at_entry_1437;
      req <= phi_stmt_1470_req_0 & phi_stmt_1470_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1470",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1470_ack_0,
          idata => idata,
          odata => input_dim0x_x1_1470,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1470
    -- flow-through select operator MUX_1579_inst
    add94_1580 <= type_cast_1577_wire_constant when (cmp_1567(0) /=  '0') else call13_1322;
    -- flow-through select operator MUX_1597_inst
    input_dim2x_x0_1598 <= add87_1582_delayed_1_0_1591 when (cmp_1567(0) /=  '0') else type_cast_1596_wire_constant;
    -- flow-through select operator MUX_1675_inst
    MUX_1675_wire <= type_cast_1645_1645_delayed_2_0_1666 when (whilex_xbody_ifx_xend122_taken_1628(0) /=  '0') else type_cast_1674_wire_constant;
    -- flow-through select operator MUX_1676_inst
    add_dest_dim0x_x0_1677 <= type_cast_1670_wire when (ifx_xthen103_ifx_xend122_taken_1662(0) /=  '0') else MUX_1675_wire;
    -- flow-through select operator MUX_1690_inst
    MUX_1690_wire <= type_cast_1657_1657_delayed_1_0_1681 when (whilex_xbody_ifx_xend122_taken_1628(0) /=  '0') else type_cast_1689_wire_constant;
    -- flow-through select operator MUX_1691_inst
    add_dest_dim1x_x2_1692 <= type_cast_1685_wire when (ifx_xthen103_ifx_xend122_taken_1662(0) /=  '0') else MUX_1690_wire;
    -- flow-through select operator MUX_1703_inst
    MUX_1703_wire <= type_cast_1700_wire when (whilex_xbody_ifx_xend122_taken_1628(0) /=  '0') else type_cast_1702_wire_constant;
    -- flow-through select operator MUX_1704_inst
    input_dim1x_x2_1705 <= type_cast_1697_wire_constant when (ifx_xthen103_ifx_xend122_taken_1662(0) /=  '0') else MUX_1703_wire;
    -- flow-through select operator MUX_1718_inst
    MUX_1718_wire <= type_cast_1682_1682_delayed_2_0_1709 when (whilex_xbody_ifx_xend122_taken_1628(0) /=  '0') else type_cast_1717_wire_constant;
    -- flow-through select operator MUX_1719_inst
    input_dim0x_x0_1720 <= type_cast_1713_wire when (ifx_xthen103_ifx_xend122_taken_1662(0) /=  '0') else MUX_1718_wire;
    W_add87_1582_delayed_1_0_1589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add87_1582_delayed_1_0_1589_inst_req_0;
      W_add87_1582_delayed_1_0_1589_inst_ack_0<= wack(0);
      rreq(0) <= W_add87_1582_delayed_1_0_1589_inst_req_1;
      W_add87_1582_delayed_1_0_1589_inst_ack_1<= rack(0);
      W_add87_1582_delayed_1_0_1589_inst : InterlockBuffer generic map ( -- 
        name => "W_add87_1582_delayed_1_0_1589_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add87_1573,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add87_1582_delayed_1_0_1591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_req_0;
      W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_ack_0<= wack(0);
      rreq(0) <= W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_req_1;
      W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst_ack_1<= rack(0);
      W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst : InterlockBuffer generic map ( -- 
        name => "W_add_dest_dim0x_x1_1626_delayed_2_0_1642_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0x_x1_1450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim0x_x1_1626_delayed_2_0_1644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_req_0;
      W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_ack_0<= wack(0);
      rreq(0) <= W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_req_1;
      W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst_ack_1<= rack(0);
      W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst : InterlockBuffer generic map ( -- 
        name => "W_add_dest_dim1x_x0_1632_delayed_1_0_1651_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1x_x0_1588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1x_x0_1632_delayed_1_0_1653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_req_0;
      W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_ack_0<= wack(0);
      rreq(0) <= W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_req_1;
      W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst_ack_1<= rack(0);
      W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst : InterlockBuffer generic map ( -- 
        name => "W_add_dest_dim1x_x1_1577_delayed_1_0_1581_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1x_x1_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1x_x1_1577_delayed_1_0_1583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx72_1547_delayed_6_0_1547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx72_1547_delayed_6_0_1547_inst_req_0;
      W_arrayidx72_1547_delayed_6_0_1547_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx72_1547_delayed_6_0_1547_inst_req_1;
      W_arrayidx72_1547_delayed_6_0_1547_inst_ack_1<= rack(0);
      W_arrayidx72_1547_delayed_6_0_1547_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx72_1547_delayed_6_0_1547_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx72_1546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx72_1547_delayed_6_0_1549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xend122_whilex_xend_taken_1736_inst
    process(cmp129_1729) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp129_1729(0 downto 0);
      ifx_xend122_whilex_xend_taken_1738 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen103_exec_guard_1629_inst
    process(whilex_xbody_ifx_xthen103_taken_1624) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xthen103_taken_1624(0 downto 0);
      ifx_xthen103_exec_guard_1631 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen103_ifx_xend122_taken_1660_inst
    process(ifx_xthen103_exec_guard_1631) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen103_exec_guard_1631(0 downto 0);
      ifx_xthen103_ifx_xend122_taken_1662 <= tmp_var; -- 
    end process;
    W_input_dim0x_x1_1619_delayed_2_0_1632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim0x_x1_1619_delayed_2_0_1632_inst_req_0;
      W_input_dim0x_x1_1619_delayed_2_0_1632_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim0x_x1_1619_delayed_2_0_1632_inst_req_1;
      W_input_dim0x_x1_1619_delayed_2_0_1632_inst_ack_1<= rack(0);
      W_input_dim0x_x1_1619_delayed_2_0_1632_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim0x_x1_1619_delayed_2_0_1632_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_1470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_1619_delayed_2_0_1634,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim1x_x1_1599_delayed_2_0_1609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim1x_x1_1599_delayed_2_0_1609_inst_req_0;
      W_input_dim1x_x1_1599_delayed_2_0_1609_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim1x_x1_1599_delayed_2_0_1609_inst_req_1;
      W_input_dim1x_x1_1599_delayed_2_0_1609_inst_ack_1<= rack(0);
      W_input_dim1x_x1_1599_delayed_2_0_1609_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim1x_x1_1599_delayed_2_0_1609_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim1x_x1_1599_delayed_2_0_1611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_ifx_xthen103_taken_1622_inst
    process(cmp101_1621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp101_1621(0 downto 0);
      whilex_xbody_ifx_xthen103_taken_1624 <= tmp_var; -- 
    end process;
    add_dest_dim0x_x1_at_entry_1419_1454_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim0x_x1_at_entry_1419_1454_buf_req_0;
      add_dest_dim0x_x1_at_entry_1419_1454_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim0x_x1_at_entry_1419_1454_buf_req_1;
      add_dest_dim0x_x1_at_entry_1419_1454_buf_ack_1<= rack(0);
      add_dest_dim0x_x1_at_entry_1419_1454_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim0x_x1_at_entry_1419_1454_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0x_x1_at_entry_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim0x_x1_at_entry_1419_1454_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim1x_x1_at_entry_1423_1459_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim1x_x1_at_entry_1423_1459_buf_req_0;
      add_dest_dim1x_x1_at_entry_1423_1459_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim1x_x1_at_entry_1423_1459_buf_req_1;
      add_dest_dim1x_x1_at_entry_1423_1459_buf_ack_1<= rack(0);
      add_dest_dim1x_x1_at_entry_1423_1459_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim1x_x1_at_entry_1423_1459_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1x_x1_at_entry_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1x_x1_at_entry_1423_1459_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1522_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1522_final_reg_req_0;
      addr_of_1522_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1522_final_reg_req_1;
      addr_of_1522_final_reg_ack_1<= rack(0);
      addr_of_1522_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1522_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1521_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx68_1523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1545_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1545_final_reg_req_0;
      addr_of_1545_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1545_final_reg_req_1;
      addr_of_1545_final_reg_ack_1<= rack(0);
      addr_of_1545_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1545_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1544_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx72_1546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1331_inst_req_0;
      type_cast_1331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1331_inst_req_1;
      type_cast_1331_inst_ack_1<= rack(0);
      type_cast_1331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1344_inst_req_0;
      type_cast_1344_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1344_inst_req_1;
      type_cast_1344_inst_ack_1<= rack(0);
      type_cast_1344_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1344_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1345,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1379_inst_req_0;
      type_cast_1379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1379_inst_req_1;
      type_cast_1379_inst_ack_1<= rack(0);
      type_cast_1379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1379_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1359,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1380,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1383_inst_req_0;
      type_cast_1383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1383_inst_req_1;
      type_cast_1383_inst_ack_1<= rack(0);
      type_cast_1383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1395_inst_req_0;
      type_cast_1395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1395_inst_req_1;
      type_cast_1395_inst_ack_1<= rack(0);
      type_cast_1395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1394_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1404_inst_req_0;
      type_cast_1404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1404_inst_req_1;
      type_cast_1404_inst_ack_1<= rack(0);
      type_cast_1404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_1405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1422_inst_req_0;
      type_cast_1422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1422_inst_req_1;
      type_cast_1422_inst_ack_1<= rack(0);
      type_cast_1422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1371,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1422_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1426_inst_req_0;
      type_cast_1426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1426_inst_req_1;
      type_cast_1426_inst_ack_1<= rack(0);
      type_cast_1426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub45_1376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1426_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1449_inst_req_0;
      type_cast_1449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1449_inst_req_1;
      type_cast_1449_inst_ack_1<= rack(0);
      type_cast_1449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1449_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1449_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1453_inst_req_0;
      type_cast_1453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1453_inst_req_1;
      type_cast_1453_inst_ack_1<= rack(0);
      type_cast_1453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1453_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0x_x0_1677,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1453_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1458_inst_req_0;
      type_cast_1458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1458_inst_req_1;
      type_cast_1458_inst_ack_1<= rack(0);
      type_cast_1458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1458_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1x_x2_1692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1458_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1463_inst_req_0;
      type_cast_1463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1463_inst_req_1;
      type_cast_1463_inst_ack_1<= rack(0);
      type_cast_1463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1463_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0_1598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1463_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1468_inst_req_0;
      type_cast_1468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1468_inst_req_1;
      type_cast_1468_inst_ack_1<= rack(0);
      type_cast_1468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1468_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1468_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1473_inst_req_0;
      type_cast_1473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1473_inst_req_1;
      type_cast_1473_inst_ack_1<= rack(0);
      type_cast_1473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1473_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1720,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1473_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1483_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1483_inst_req_0;
      type_cast_1483_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1483_inst_req_1;
      type_cast_1483_inst_ack_1<= rack(0);
      type_cast_1483_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1483_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1487_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1487_inst_req_0;
      type_cast_1487_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1487_inst_req_1;
      type_cast_1487_inst_ack_1<= rack(0);
      type_cast_1487_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1487_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1x_x1_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_1488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1491_inst_req_0;
      type_cast_1491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1491_inst_req_1;
      type_cast_1491_inst_ack_1<= rack(0);
      type_cast_1491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0x_x1_1450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_1492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1515_inst_req_0;
      type_cast_1515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1515_inst_req_1;
      type_cast_1515_inst_ack_1<= rack(0);
      type_cast_1515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_src_0x_x0_1480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1556_inst_req_0;
      type_cast_1556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1556_inst_req_1;
      type_cast_1556_inst_ack_1<= rack(0);
      type_cast_1556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1556_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1560_inst_req_0;
      type_cast_1560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1560_inst_req_1;
      type_cast_1560_inst_ack_1<= rack(0);
      type_cast_1560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1560_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv83_1396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1559_1559_delayed_2_0_1561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1564_inst
    process(conv81_1557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv81_1557(31 downto 0);
      type_cast_1564_wire <= tmp_var; -- 
    end process;
    type_cast_1601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1601_inst_req_0;
      type_cast_1601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1601_inst_req_1;
      type_cast_1601_inst_ack_1<= rack(0);
      type_cast_1601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1601_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_1567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_18_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1665_inst_req_0;
      type_cast_1665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1665_inst_req_1;
      type_cast_1665_inst_ack_1<= rack(0);
      type_cast_1665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1665_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0x_x1_1450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1645_1645_delayed_2_0_1666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1670_inst
    process(add110_1650) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add110_1650(15 downto 0);
      type_cast_1670_wire <= tmp_var; -- 
    end process;
    type_cast_1680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1680_inst_req_0;
      type_cast_1680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1680_inst_req_1;
      type_cast_1680_inst_ack_1<= rack(0);
      type_cast_1680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1680_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1x_x0_1588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1657_1657_delayed_1_0_1681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1685_inst
    process(sub120_1659) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sub120_1659(15 downto 0);
      type_cast_1685_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1700_inst
    process(input_dim1x_x0_1616) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := input_dim1x_x0_1616(15 downto 0);
      type_cast_1700_wire <= tmp_var; -- 
    end process;
    type_cast_1708_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1708_inst_req_0;
      type_cast_1708_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1708_inst_req_1;
      type_cast_1708_inst_ack_1<= rack(0);
      type_cast_1708_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1708_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_1470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1682_1682_delayed_2_0_1709,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1713_inst
    process(inc105_1641) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc105_1641(15 downto 0);
      type_cast_1713_wire <= tmp_var; -- 
    end process;
    type_cast_1723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1723_inst_req_0;
      type_cast_1723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1723_inst_req_1;
      type_cast_1723_inst_ack_1<= rack(0);
      type_cast_1723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1720,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv124_1724,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1521_index_1_rename
    process(R_idxprom_1520_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1520_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1520_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1521_index_1_resize
    process(idxprom_1516) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1516;
      ov := iv(13 downto 0);
      R_idxprom_1520_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1521_root_address_inst
    process(array_obj_ref_1521_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1521_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1521_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1544_index_1_rename
    process(R_idxprom71_1543_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom71_1543_resized;
      ov(13 downto 0) := iv;
      R_idxprom71_1543_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1544_index_1_resize
    process(idxprom71_1539) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom71_1539;
      ov := iv(13 downto 0);
      R_idxprom71_1543_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1544_root_address_inst
    process(array_obj_ref_1544_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1544_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1544_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_addr_0
    process(ptr_deref_1526_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1526_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1526_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_base_resize
    process(arrayidx68_1523) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx68_1523;
      ov := iv(13 downto 0);
      ptr_deref_1526_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_gather_scatter
    process(ptr_deref_1526_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1526_data_0;
      ov(63 downto 0) := iv;
      tmp69_1527 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_root_address_inst
    process(ptr_deref_1526_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1526_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1526_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_addr_0
    process(ptr_deref_1551_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1551_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1551_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_base_resize
    process(arrayidx72_1547_delayed_6_0_1549) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx72_1547_delayed_6_0_1549;
      ov := iv(13 downto 0);
      ptr_deref_1551_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_gather_scatter
    process(tmp69_1527) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp69_1527;
      ov(63 downto 0) := iv;
      ptr_deref_1551_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_root_address_inst
    process(ptr_deref_1551_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1551_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1551_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_1443_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1741_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1443_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1443_branch_req_0,
          ack0 => do_while_stmt_1443_branch_ack_0,
          ack1 => do_while_stmt_1443_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1742_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ifx_xend122_whilex_xend_taken_1738;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1742_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1742_branch_req_0,
          ack0 => if_stmt_1742_branch_ack_0,
          ack1 => if_stmt_1742_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1365_inst
    process(call14_1325) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call14_1325, type_cast_1364_wire_constant, tmp_var);
      add30_1366 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1389_inst
    process(call3_1307) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call3_1307, type_cast_1388_wire_constant, tmp_var);
      sub77_1390 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1572_inst
    process(input_dim2x_x1_1460) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1460, type_cast_1571_wire_constant, tmp_var);
      add87_1573 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1587_inst
    process(add94_1580, add_dest_dim1x_x1_1577_delayed_1_0_1583) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add94_1580, add_dest_dim1x_x1_1577_delayed_1_0_1583, tmp_var);
      add_dest_dim1x_x0_1588 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1615_inst
    process(inc_1608, input_dim1x_x1_1599_delayed_2_0_1611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc_1608, input_dim1x_x1_1599_delayed_2_0_1611, tmp_var);
      input_dim1x_x0_1616 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1640_inst
    process(input_dim0x_x1_1619_delayed_2_0_1634) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x1_1619_delayed_2_0_1634, type_cast_1639_wire_constant, tmp_var);
      inc105_1641 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1649_inst
    process(add_dest_dim0x_x1_1626_delayed_2_0_1644, call13_1322) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim0x_x1_1626_delayed_2_0_1644, call13_1322, tmp_var);
      add110_1650 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1479_inst
    process(add_1350, indvar_1445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1350, indvar_1445, tmp_var);
      add_src_0x_x0_1480 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1734_inst
    process(indvar_1445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1445, type_cast_1733_wire_constant, tmp_var);
      indvarx_xnext_1735 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1501_inst
    process(conv58_1488, mul_1497) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv58_1488, mul_1497, tmp_var);
      add64_1502 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1511_inst
    process(mul65_1507, conv53_1484) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul65_1507, conv53_1484, tmp_var);
      add66_1512 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1538_inst
    process(shr_1533) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr_1533, type_cast_1537_wire_constant, tmp_var);
      idxprom71_1539 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1620_inst
    process(input_dim1x_x0_1616, call1_1304) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1x_x0_1616, call1_1304, tmp_var);
      cmp101_1621 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1728_inst
    process(conv124_1724, shr128142_1411) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv124_1724, shr128142_1411, tmp_var);
      cmp129_1729 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1410_inst
    process(conv127_1405) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv127_1405, type_cast_1409_wire_constant, tmp_var);
      shr128142_1411 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1532_inst
    process(add66_1512) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add66_1512, type_cast_1531_wire_constant, tmp_var);
      shr_1533 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1400_inst
    process(call13_1322, call1_1304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1322, call1_1304, tmp_var);
      mul117_1401 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1496_inst
    process(conv63_1492, conv61_1384) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_1492, conv61_1384, tmp_var);
      mul_1497 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1506_inst
    process(add64_1502, conv56_1380) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add64_1502, conv56_1380, tmp_var);
      mul65_1507 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1627_inst
    process(cmp101_1621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp101_1621, tmp_var);
      whilex_xbody_ifx_xend122_taken_1628 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1741_inst
    process(cmp129_1729) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp129_1729, tmp_var);
      NOT_u1_u1_1741_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u32_u32_1349_inst
    process(shl_1338, conv17_1345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1338, conv17_1345, tmp_var);
      add_1350 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1337_inst
    process(conv_1332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1332, type_cast_1336_wire_constant, tmp_var);
      shl_1338 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1566_inst
    process(type_cast_1564_wire, type_cast_1559_1559_delayed_2_0_1561) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1564_wire, type_cast_1559_1559_delayed_2_0_1561, tmp_var);
      cmp_1567 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1370_inst
    process(call7_1313, add30_1366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(call7_1313, add30_1366, tmp_var);
      sub_1371 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1375_inst
    process(call9_1316, add30_1366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(call9_1316, add30_1366, tmp_var);
      sub45_1376 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1658_inst
    process(add_dest_dim1x_x0_1632_delayed_1_0_1653, mul117_1401) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add_dest_dim1x_x0_1632_delayed_1_0_1653, mul117_1401, tmp_var);
      sub120_1659 <= tmp_var; --
    end process;
    -- binary operator XOR_u16_u16_1607_inst
    process(iNsTr_18_1602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntXor_proc(iNsTr_18_1602, type_cast_1606_wire_constant, tmp_var);
      inc_1608 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1521_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1520_scaled;
      array_obj_ref_1521_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1521_index_offset_req_0;
      array_obj_ref_1521_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1521_index_offset_req_1;
      array_obj_ref_1521_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1544_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom71_1543_scaled;
      array_obj_ref_1544_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1544_index_offset_req_0;
      array_obj_ref_1544_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1544_index_offset_req_1;
      array_obj_ref_1544_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1394_inst
    process(sub77_1390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", sub77_1390, tmp_var);
      type_cast_1394_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1526_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1526_load_0_req_0;
      ptr_deref_1526_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1526_load_0_req_1;
      ptr_deref_1526_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1526_word_address_0;
      ptr_deref_1526_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1551_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1551_store_0_req_0;
      ptr_deref_1551_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1551_store_0_req_1;
      ptr_deref_1551_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1551_word_address_0;
      data_in <= ptr_deref_1551_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1300_inst RPIPE_Block0_start_1303_inst RPIPE_Block0_start_1306_inst RPIPE_Block0_start_1309_inst RPIPE_Block0_start_1312_inst RPIPE_Block0_start_1315_inst RPIPE_Block0_start_1318_inst RPIPE_Block0_start_1321_inst RPIPE_Block0_start_1324_inst RPIPE_Block0_start_1327_inst RPIPE_Block0_start_1340_inst RPIPE_Block0_start_1352_inst RPIPE_Block0_start_1355_inst RPIPE_Block0_start_1358_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1300_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1303_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1306_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1309_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1312_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1315_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1318_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1321_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1324_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1327_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1340_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1352_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1355_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1358_inst_req_0;
      RPIPE_Block0_start_1300_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1303_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1306_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1309_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1312_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1315_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1318_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1321_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1324_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1327_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1340_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1352_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1355_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1358_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1300_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1303_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1306_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1309_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1312_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1315_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1318_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1321_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1324_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1327_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1340_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1352_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1355_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1358_inst_req_1;
      RPIPE_Block0_start_1300_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1303_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1306_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1309_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1312_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1315_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1318_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1321_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1324_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1327_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1340_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1352_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1355_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1358_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_1301 <= data_out(223 downto 208);
      call1_1304 <= data_out(207 downto 192);
      call3_1307 <= data_out(191 downto 176);
      call5_1310 <= data_out(175 downto 160);
      call7_1313 <= data_out(159 downto 144);
      call9_1316 <= data_out(143 downto 128);
      call11_1319 <= data_out(127 downto 112);
      call13_1322 <= data_out(111 downto 96);
      call14_1325 <= data_out(95 downto 80);
      call15_1328 <= data_out(79 downto 64);
      call16_1341 <= data_out(63 downto 48);
      call18_1353 <= data_out(47 downto 32);
      call20_1356 <= data_out(31 downto 16);
      call22_1359 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1748_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1748_inst_req_0;
      WPIPE_Block0_done_1748_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1748_inst_req_1;
      WPIPE_Block0_done_1748_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1750_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_23_inst_req_0 : boolean;
  signal WPIPE_timer_req_23_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_28_inst_req_0 : boolean;
  signal RPIPE_timer_resp_28_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_28_inst_req_1 : boolean;
  signal RPIPE_timer_resp_28_inst_ack_1 : boolean;
  signal WPIPE_timer_req_23_inst_req_1 : boolean;
  signal WPIPE_timer_req_23_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Sample/req
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Sample/rr
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/$entry
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_sample_start_
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_sample_start_
      -- CP-element group 0: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Sample/$entry
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_28_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_23_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Sample/ack
      -- CP-element group 1: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_sample_completed_
      -- CP-element group 1: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_update_start_
      -- CP-element group 1: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Update/$entry
      -- CP-element group 1: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_23_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_23_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_update_completed_
      -- CP-element group 2: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Update/$exit
      -- CP-element group 2: 	 assign_stmt_26_to_assign_stmt_29/WPIPE_timer_req_23_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_23_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Sample/ra
      -- CP-element group 3: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Update/$entry
      -- CP-element group 3: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Update/cr
      -- CP-element group 3: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_sample_completed_
      -- CP-element group 3: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_update_start_
      -- CP-element group 3: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Sample/$exit
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_28_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_28_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Update/$exit
      -- CP-element group 4: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_Update/ca
      -- CP-element group 4: 	 assign_stmt_26_to_assign_stmt_29/RPIPE_timer_resp_28_update_completed_
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_28_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_26_to_assign_stmt_29/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(2) & timer_CP_0_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_25_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_25_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_28_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_28_inst_req_0;
      RPIPE_timer_resp_28_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_28_inst_req_1;
      RPIPE_timer_resp_28_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_23_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_23_inst_req_0;
      WPIPE_timer_req_23_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_23_inst_req_1;
      WPIPE_timer_req_23_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_25_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_4253_start: Boolean;
  signal timerDaemon_CP_4253_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1766_branch_req_0 : boolean;
  signal phi_stmt_1768_req_0 : boolean;
  signal phi_stmt_1768_req_1 : boolean;
  signal phi_stmt_1768_ack_0 : boolean;
  signal nCOUNTER_1781_1770_buf_req_0 : boolean;
  signal nCOUNTER_1781_1770_buf_ack_0 : boolean;
  signal nCOUNTER_1781_1770_buf_req_1 : boolean;
  signal nCOUNTER_1781_1770_buf_ack_1 : boolean;
  signal RPIPE_timer_req_1775_inst_req_0 : boolean;
  signal RPIPE_timer_req_1775_inst_ack_0 : boolean;
  signal RPIPE_timer_req_1775_inst_req_1 : boolean;
  signal RPIPE_timer_req_1775_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_1783_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1783_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_1783_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1783_inst_ack_1 : boolean;
  signal do_while_stmt_1766_branch_ack_0 : boolean;
  signal do_while_stmt_1766_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_4253_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4253_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_4253_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4253_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_4253: Block -- control-path 
    signal timerDaemon_CP_4253_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_4253_elements(0) <= timerDaemon_CP_4253_start;
    timerDaemon_CP_4253_symbol <= timerDaemon_CP_4253_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1765/$entry
      -- CP-element group 0: 	 branch_block_stmt_1765/branch_block_stmt_1765__entry__
      -- CP-element group 0: 	 branch_block_stmt_1765/do_while_stmt_1766__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1765/$exit
      -- CP-element group 1: 	 branch_block_stmt_1765/branch_block_stmt_1765__exit__
      -- CP-element group 1: 	 branch_block_stmt_1765/do_while_stmt_1766__exit__
      -- 
    timerDaemon_CP_4253_elements(1) <= timerDaemon_CP_4253_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1765/do_while_stmt_1766/$entry
      -- CP-element group 2: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766__entry__
      -- 
    timerDaemon_CP_4253_elements(2) <= timerDaemon_CP_4253_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766__exit__
      -- 
    -- Element group timerDaemon_CP_4253_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_back
      -- 
    -- Element group timerDaemon_CP_4253_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1765/do_while_stmt_1766/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_taken/$entry
      -- 
    timerDaemon_CP_4253_elements(5) <= timerDaemon_CP_4253_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_body_done
      -- 
    timerDaemon_CP_4253_elements(6) <= timerDaemon_CP_4253_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_4253_elements(7) <= timerDaemon_CP_4253_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_4253_elements(8) <= timerDaemon_CP_4253_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1773_sample_start_
      -- 
    -- Element group timerDaemon_CP_4253_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/condition_evaluated
      -- 
    condition_evaluated_4277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(10), ack => do_while_stmt_1766_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(40) & timerDaemon_CP_4253_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(9) & timerDaemon_CP_4253_elements(15) & timerDaemon_CP_4253_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1773_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(35) & timerDaemon_CP_4253_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(32) & timerDaemon_CP_4253_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(36) & timerDaemon_CP_4253_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(9) & timerDaemon_CP_4253_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(9) & timerDaemon_CP_4253_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_4253_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_4253_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_loopback_trigger
      -- 
    timerDaemon_CP_4253_elements(19) <= timerDaemon_CP_4253_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_loopback_sample_req_ps
      -- 
    phi_stmt_1768_loopback_sample_req_4292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1768_loopback_sample_req_4292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(20), ack => phi_stmt_1768_req_0); -- 
    -- Element group timerDaemon_CP_4253_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_entry_trigger
      -- 
    timerDaemon_CP_4253_elements(21) <= timerDaemon_CP_4253_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_entry_sample_req_ps
      -- 
    phi_stmt_1768_entry_sample_req_4295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1768_entry_sample_req_4295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(22), ack => phi_stmt_1768_req_1); -- 
    -- Element group timerDaemon_CP_4253_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1768_phi_mux_ack_ps
      -- 
    phi_stmt_1768_phi_mux_ack_4298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1768_ack_0, ack => timerDaemon_CP_4253_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Sample/req
      -- 
    req_4311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(24), ack => nCOUNTER_1781_1770_buf_req_0); -- 
    -- Element group timerDaemon_CP_4253_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Update/req
      -- 
    req_4316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(25), ack => nCOUNTER_1781_1770_buf_req_1); -- 
    -- Element group timerDaemon_CP_4253_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Sample/ack
      -- 
    ack_4312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1781_1770_buf_ack_0, ack => timerDaemon_CP_4253_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/R_nCOUNTER_1770_Update/ack
      -- 
    ack_4317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1781_1770_buf_ack_1, ack => timerDaemon_CP_4253_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_sample_completed_
      -- 
    -- Element group timerDaemon_CP_4253_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_update_start_
      -- 
    -- Element group timerDaemon_CP_4253_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_update_completed__ps
      -- 
    timerDaemon_CP_4253_elements(30) <= timerDaemon_CP_4253_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/type_cast_1772_update_completed_
      -- 
    -- Element group timerDaemon_CP_4253_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => timerDaemon_CP_4253_elements(29), ack => timerDaemon_CP_4253_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1773_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(9) & timerDaemon_CP_4253_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Sample/rr
      -- 
    rr_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(33), ack => RPIPE_timer_req_1775_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(11) & timerDaemon_CP_4253_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Update/cr
      -- 
    cr_4343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(34), ack => RPIPE_timer_req_1775_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(35) & timerDaemon_CP_4253_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Sample/ra
      -- 
    ra_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1775_inst_ack_0, ack => timerDaemon_CP_4253_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/phi_stmt_1773_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/RPIPE_timer_req_1775_Update/ca
      -- 
    ca_4344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1775_inst_ack_1, ack => timerDaemon_CP_4253_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Sample/req
      -- 
    req_4352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(37), ack => WPIPE_timer_resp_1783_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(36) & timerDaemon_CP_4253_elements(18) & timerDaemon_CP_4253_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Update/req
      -- 
    ack_4353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1783_inst_ack_0, ack => timerDaemon_CP_4253_elements(38)); -- 
    req_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4253_elements(38), ack => WPIPE_timer_resp_1783_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/WPIPE_timer_resp_1783_Update/ack
      -- 
    ack_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1783_inst_ack_1, ack => timerDaemon_CP_4253_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_4253_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_4253_elements(9), ack => timerDaemon_CP_4253_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1765/do_while_stmt_1766/do_while_stmt_1766_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4253_elements(39) & timerDaemon_CP_4253_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4253_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_exit/ack
      -- 
    ack_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1766_branch_ack_0, ack => timerDaemon_CP_4253_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1765/do_while_stmt_1766/loop_taken/ack
      -- 
    ack_4367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1766_branch_ack_1, ack => timerDaemon_CP_4253_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1765/do_while_stmt_1766/$exit
      -- 
    timerDaemon_CP_4253_elements(44) <= timerDaemon_CP_4253_elements(3);
    timerDaemon_do_while_stmt_1766_terminator_4368: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1766_terminator_4368", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_4253_elements(6),loop_continue => timerDaemon_CP_4253_elements(43),loop_terminate => timerDaemon_CP_4253_elements(42),loop_back => timerDaemon_CP_4253_elements(4),loop_exit => timerDaemon_CP_4253_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1768_phi_seq_4326_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_4253_elements(19);
      timerDaemon_CP_4253_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_4253_elements(26);
      timerDaemon_CP_4253_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_4253_elements(27);
      timerDaemon_CP_4253_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_4253_elements(21);
      timerDaemon_CP_4253_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_4253_elements(28);
      timerDaemon_CP_4253_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_4253_elements(30);
      timerDaemon_CP_4253_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1768_phi_seq_4326 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1768_phi_seq_4326") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_4253_elements(11), 
          phi_sample_ack => timerDaemon_CP_4253_elements(17), 
          phi_update_req => timerDaemon_CP_4253_elements(13), 
          phi_update_ack => timerDaemon_CP_4253_elements(18), 
          phi_mux_ack => timerDaemon_CP_4253_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4278_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_4253_elements(7);
        preds(1)  <= timerDaemon_CP_4253_elements(8);
        entry_tmerge_4278 : transition_merge -- 
          generic map(name => " entry_tmerge_4278")
          port map (preds => preds, symbol_out => timerDaemon_CP_4253_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1768 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1775_wire : std_logic_vector(0 downto 0);
    signal konst_1779_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1787_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1781 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1781_1770_buffered : std_logic_vector(63 downto 0);
    signal req_1773 : std_logic_vector(0 downto 0);
    signal type_cast_1772_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1779_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1787_wire_constant <= "1";
    type_cast_1772_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1768: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nCOUNTER_1781_1770_buffered & type_cast_1772_wire_constant;
      req <= phi_stmt_1768_req_0 & phi_stmt_1768_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1768",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1768_ack_0,
          idata => idata,
          odata => COUNTER_1768,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1768
    nCOUNTER_1781_1770_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1781_1770_buf_req_0;
      nCOUNTER_1781_1770_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1781_1770_buf_req_1;
      nCOUNTER_1781_1770_buf_ack_1<= rack(0);
      nCOUNTER_1781_1770_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1781_1770_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1781_1770_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1773
    process(RPIPE_timer_req_1775_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1775_wire(0 downto 0);
      req_1773 <= tmp_var; -- 
    end process;
    do_while_stmt_1766_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1787_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1766_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1766_branch_req_0,
          ack0 => do_while_stmt_1766_branch_ack_0,
          ack1 => do_while_stmt_1766_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1780_inst
    process(COUNTER_1768) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1768, konst_1779_wire_constant, tmp_var);
      nCOUNTER_1781 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1775_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1775_inst_req_0;
      RPIPE_timer_req_1775_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1775_inst_req_1;
      RPIPE_timer_req_1775_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1775_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1783_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1783_inst_req_0;
      WPIPE_timer_resp_1783_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1783_inst_req_1;
      WPIPE_timer_resp_1783_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1773(0);
      data_in <= COUNTER_1768;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(27 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(35 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(10 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(27 downto 14),
      memory_space_2_sr_data => memory_space_2_sr_data(127 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(35 downto 18),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 2,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
